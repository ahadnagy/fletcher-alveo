-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.Array_pkg.all;
use work.mmio_pkg.all;

entity Kernel_Nucleus is
  generic (
    INDEX_WIDTH                        : integer := 32;
    TAG_WIDTH                          : integer := 1;
    REMATCH000_IN_BUS_ADDR_WIDTH       : integer := 64;
    REMATCH001_IN_BUS_ADDR_WIDTH       : integer := 64;
    REMATCH002_IN_BUS_ADDR_WIDTH       : integer := 64;
    REMATCH003_IN_BUS_ADDR_WIDTH       : integer := 64;
    REMATCH004_IN_BUS_ADDR_WIDTH       : integer := 64;
    REMATCH005_IN_BUS_ADDR_WIDTH       : integer := 64;
    REMATCH006_IN_BUS_ADDR_WIDTH       : integer := 64;
    REMATCH007_IN_BUS_ADDR_WIDTH       : integer := 64;
    REMATCH008_IN_BUS_ADDR_WIDTH       : integer := 64;
    REMATCH009_IN_BUS_ADDR_WIDTH       : integer := 64;
    REMATCH010_IN_BUS_ADDR_WIDTH       : integer := 64;
    REMATCH011_IN_BUS_ADDR_WIDTH       : integer := 64;
    REMATCH012_IN_BUS_ADDR_WIDTH       : integer := 64;
    REMATCH013_IN_BUS_ADDR_WIDTH       : integer := 64;
    REMATCH014_IN_BUS_ADDR_WIDTH       : integer := 64;
    REMATCH015_IN_BUS_ADDR_WIDTH       : integer := 64;
    REMATCH000_TAXI_OUT_BUS_ADDR_WIDTH : integer := 64;
    REMATCH001_TAXI_OUT_BUS_ADDR_WIDTH : integer := 64;
    REMATCH002_TAXI_OUT_BUS_ADDR_WIDTH : integer := 64;
    REMATCH003_TAXI_OUT_BUS_ADDR_WIDTH : integer := 64;
    REMATCH004_TAXI_OUT_BUS_ADDR_WIDTH : integer := 64;
    REMATCH005_TAXI_OUT_BUS_ADDR_WIDTH : integer := 64;
    REMATCH006_TAXI_OUT_BUS_ADDR_WIDTH : integer := 64;
    REMATCH007_TAXI_OUT_BUS_ADDR_WIDTH : integer := 64;
    REMATCH008_TAXI_OUT_BUS_ADDR_WIDTH : integer := 64;
    REMATCH009_TAXI_OUT_BUS_ADDR_WIDTH : integer := 64;
    REMATCH010_TAXI_OUT_BUS_ADDR_WIDTH : integer := 64;
    REMATCH011_TAXI_OUT_BUS_ADDR_WIDTH : integer := 64;
    REMATCH012_TAXI_OUT_BUS_ADDR_WIDTH : integer := 64;
    REMATCH013_TAXI_OUT_BUS_ADDR_WIDTH : integer := 64;
    REMATCH014_TAXI_OUT_BUS_ADDR_WIDTH : integer := 64;
    REMATCH015_TAXI_OUT_BUS_ADDR_WIDTH : integer := 64
  );
  port (
    kcd_clk                          : in  std_logic;
    kcd_reset                        : in  std_logic;
    mmio_awvalid                     : in  std_logic;
    mmio_awready                     : out std_logic;
    mmio_awaddr                      : in  std_logic_vector(31 downto 0);
    mmio_wvalid                      : in  std_logic;
    mmio_wready                      : out std_logic;
    mmio_wdata                       : in  std_logic_vector(31 downto 0);
    mmio_wstrb                       : in  std_logic_vector(3 downto 0);
    mmio_bvalid                      : out std_logic;
    mmio_bready                      : in  std_logic;
    mmio_bresp                       : out std_logic_vector(1 downto 0);
    mmio_arvalid                     : in  std_logic;
    mmio_arready                     : out std_logic;
    mmio_araddr                      : in  std_logic_vector(31 downto 0);
    mmio_rvalid                      : out std_logic;
    mmio_rready                      : in  std_logic;
    mmio_rdata                       : out std_logic_vector(31 downto 0);
    mmio_rresp                       : out std_logic_vector(1 downto 0);
    rematch000_in_valid              : in  std_logic;
    rematch000_in_ready              : out std_logic;
    rematch000_in_dvalid             : in  std_logic;
    rematch000_in_last               : in  std_logic;
    rematch000_in_length             : in  std_logic_vector(31 downto 0);
    rematch000_in_count              : in  std_logic_vector(0 downto 0);
    rematch000_in_chars_valid        : in  std_logic;
    rematch000_in_chars_ready        : out std_logic;
    rematch000_in_chars_dvalid       : in  std_logic;
    rematch000_in_chars_last         : in  std_logic;
    rematch000_in_chars              : in  std_logic_vector(31 downto 0);
    rematch000_in_chars_count        : in  std_logic_vector(2 downto 0);
    rematch000_in_unl_valid          : in  std_logic;
    rematch000_in_unl_ready          : out std_logic;
    rematch000_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch000_in_cmd_valid          : out std_logic;
    rematch000_in_cmd_ready          : in  std_logic;
    rematch000_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch000_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch000_in_cmd_ctrl           : out std_logic_vector(REMATCH000_IN_BUS_ADDR_WIDTH*2-1 downto 0);
    rematch000_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch001_in_valid              : in  std_logic;
    rematch001_in_ready              : out std_logic;
    rematch001_in_dvalid             : in  std_logic;
    rematch001_in_last               : in  std_logic;
    rematch001_in_length             : in  std_logic_vector(31 downto 0);
    rematch001_in_count              : in  std_logic_vector(0 downto 0);
    rematch001_in_chars_valid        : in  std_logic;
    rematch001_in_chars_ready        : out std_logic;
    rematch001_in_chars_dvalid       : in  std_logic;
    rematch001_in_chars_last         : in  std_logic;
    rematch001_in_chars              : in  std_logic_vector(31 downto 0);
    rematch001_in_chars_count        : in  std_logic_vector(2 downto 0);
    rematch001_in_unl_valid          : in  std_logic;
    rematch001_in_unl_ready          : out std_logic;
    rematch001_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch001_in_cmd_valid          : out std_logic;
    rematch001_in_cmd_ready          : in  std_logic;
    rematch001_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch001_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch001_in_cmd_ctrl           : out std_logic_vector(REMATCH001_IN_BUS_ADDR_WIDTH*2-1 downto 0);
    rematch001_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch002_in_valid              : in  std_logic;
    rematch002_in_ready              : out std_logic;
    rematch002_in_dvalid             : in  std_logic;
    rematch002_in_last               : in  std_logic;
    rematch002_in_length             : in  std_logic_vector(31 downto 0);
    rematch002_in_count              : in  std_logic_vector(0 downto 0);
    rematch002_in_chars_valid        : in  std_logic;
    rematch002_in_chars_ready        : out std_logic;
    rematch002_in_chars_dvalid       : in  std_logic;
    rematch002_in_chars_last         : in  std_logic;
    rematch002_in_chars              : in  std_logic_vector(31 downto 0);
    rematch002_in_chars_count        : in  std_logic_vector(2 downto 0);
    rematch002_in_unl_valid          : in  std_logic;
    rematch002_in_unl_ready          : out std_logic;
    rematch002_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch002_in_cmd_valid          : out std_logic;
    rematch002_in_cmd_ready          : in  std_logic;
    rematch002_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch002_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch002_in_cmd_ctrl           : out std_logic_vector(REMATCH002_IN_BUS_ADDR_WIDTH*2-1 downto 0);
    rematch002_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch003_in_valid              : in  std_logic;
    rematch003_in_ready              : out std_logic;
    rematch003_in_dvalid             : in  std_logic;
    rematch003_in_last               : in  std_logic;
    rematch003_in_length             : in  std_logic_vector(31 downto 0);
    rematch003_in_count              : in  std_logic_vector(0 downto 0);
    rematch003_in_chars_valid        : in  std_logic;
    rematch003_in_chars_ready        : out std_logic;
    rematch003_in_chars_dvalid       : in  std_logic;
    rematch003_in_chars_last         : in  std_logic;
    rematch003_in_chars              : in  std_logic_vector(31 downto 0);
    rematch003_in_chars_count        : in  std_logic_vector(2 downto 0);
    rematch003_in_unl_valid          : in  std_logic;
    rematch003_in_unl_ready          : out std_logic;
    rematch003_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch003_in_cmd_valid          : out std_logic;
    rematch003_in_cmd_ready          : in  std_logic;
    rematch003_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch003_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch003_in_cmd_ctrl           : out std_logic_vector(REMATCH003_IN_BUS_ADDR_WIDTH*2-1 downto 0);
    rematch003_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch004_in_valid              : in  std_logic;
    rematch004_in_ready              : out std_logic;
    rematch004_in_dvalid             : in  std_logic;
    rematch004_in_last               : in  std_logic;
    rematch004_in_length             : in  std_logic_vector(31 downto 0);
    rematch004_in_count              : in  std_logic_vector(0 downto 0);
    rematch004_in_chars_valid        : in  std_logic;
    rematch004_in_chars_ready        : out std_logic;
    rematch004_in_chars_dvalid       : in  std_logic;
    rematch004_in_chars_last         : in  std_logic;
    rematch004_in_chars              : in  std_logic_vector(31 downto 0);
    rematch004_in_chars_count        : in  std_logic_vector(2 downto 0);
    rematch004_in_unl_valid          : in  std_logic;
    rematch004_in_unl_ready          : out std_logic;
    rematch004_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch004_in_cmd_valid          : out std_logic;
    rematch004_in_cmd_ready          : in  std_logic;
    rematch004_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch004_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch004_in_cmd_ctrl           : out std_logic_vector(REMATCH004_IN_BUS_ADDR_WIDTH*2-1 downto 0);
    rematch004_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch005_in_valid              : in  std_logic;
    rematch005_in_ready              : out std_logic;
    rematch005_in_dvalid             : in  std_logic;
    rematch005_in_last               : in  std_logic;
    rematch005_in_length             : in  std_logic_vector(31 downto 0);
    rematch005_in_count              : in  std_logic_vector(0 downto 0);
    rematch005_in_chars_valid        : in  std_logic;
    rematch005_in_chars_ready        : out std_logic;
    rematch005_in_chars_dvalid       : in  std_logic;
    rematch005_in_chars_last         : in  std_logic;
    rematch005_in_chars              : in  std_logic_vector(31 downto 0);
    rematch005_in_chars_count        : in  std_logic_vector(2 downto 0);
    rematch005_in_unl_valid          : in  std_logic;
    rematch005_in_unl_ready          : out std_logic;
    rematch005_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch005_in_cmd_valid          : out std_logic;
    rematch005_in_cmd_ready          : in  std_logic;
    rematch005_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch005_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch005_in_cmd_ctrl           : out std_logic_vector(REMATCH005_IN_BUS_ADDR_WIDTH*2-1 downto 0);
    rematch005_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch006_in_valid              : in  std_logic;
    rematch006_in_ready              : out std_logic;
    rematch006_in_dvalid             : in  std_logic;
    rematch006_in_last               : in  std_logic;
    rematch006_in_length             : in  std_logic_vector(31 downto 0);
    rematch006_in_count              : in  std_logic_vector(0 downto 0);
    rematch006_in_chars_valid        : in  std_logic;
    rematch006_in_chars_ready        : out std_logic;
    rematch006_in_chars_dvalid       : in  std_logic;
    rematch006_in_chars_last         : in  std_logic;
    rematch006_in_chars              : in  std_logic_vector(31 downto 0);
    rematch006_in_chars_count        : in  std_logic_vector(2 downto 0);
    rematch006_in_unl_valid          : in  std_logic;
    rematch006_in_unl_ready          : out std_logic;
    rematch006_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch006_in_cmd_valid          : out std_logic;
    rematch006_in_cmd_ready          : in  std_logic;
    rematch006_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch006_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch006_in_cmd_ctrl           : out std_logic_vector(REMATCH006_IN_BUS_ADDR_WIDTH*2-1 downto 0);
    rematch006_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch007_in_valid              : in  std_logic;
    rematch007_in_ready              : out std_logic;
    rematch007_in_dvalid             : in  std_logic;
    rematch007_in_last               : in  std_logic;
    rematch007_in_length             : in  std_logic_vector(31 downto 0);
    rematch007_in_count              : in  std_logic_vector(0 downto 0);
    rematch007_in_chars_valid        : in  std_logic;
    rematch007_in_chars_ready        : out std_logic;
    rematch007_in_chars_dvalid       : in  std_logic;
    rematch007_in_chars_last         : in  std_logic;
    rematch007_in_chars              : in  std_logic_vector(31 downto 0);
    rematch007_in_chars_count        : in  std_logic_vector(2 downto 0);
    rematch007_in_unl_valid          : in  std_logic;
    rematch007_in_unl_ready          : out std_logic;
    rematch007_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch007_in_cmd_valid          : out std_logic;
    rematch007_in_cmd_ready          : in  std_logic;
    rematch007_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch007_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch007_in_cmd_ctrl           : out std_logic_vector(REMATCH007_IN_BUS_ADDR_WIDTH*2-1 downto 0);
    rematch007_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch008_in_valid              : in  std_logic;
    rematch008_in_ready              : out std_logic;
    rematch008_in_dvalid             : in  std_logic;
    rematch008_in_last               : in  std_logic;
    rematch008_in_length             : in  std_logic_vector(31 downto 0);
    rematch008_in_count              : in  std_logic_vector(0 downto 0);
    rematch008_in_chars_valid        : in  std_logic;
    rematch008_in_chars_ready        : out std_logic;
    rematch008_in_chars_dvalid       : in  std_logic;
    rematch008_in_chars_last         : in  std_logic;
    rematch008_in_chars              : in  std_logic_vector(31 downto 0);
    rematch008_in_chars_count        : in  std_logic_vector(2 downto 0);
    rematch008_in_unl_valid          : in  std_logic;
    rematch008_in_unl_ready          : out std_logic;
    rematch008_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch008_in_cmd_valid          : out std_logic;
    rematch008_in_cmd_ready          : in  std_logic;
    rematch008_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch008_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch008_in_cmd_ctrl           : out std_logic_vector(REMATCH008_IN_BUS_ADDR_WIDTH*2-1 downto 0);
    rematch008_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch009_in_valid              : in  std_logic;
    rematch009_in_ready              : out std_logic;
    rematch009_in_dvalid             : in  std_logic;
    rematch009_in_last               : in  std_logic;
    rematch009_in_length             : in  std_logic_vector(31 downto 0);
    rematch009_in_count              : in  std_logic_vector(0 downto 0);
    rematch009_in_chars_valid        : in  std_logic;
    rematch009_in_chars_ready        : out std_logic;
    rematch009_in_chars_dvalid       : in  std_logic;
    rematch009_in_chars_last         : in  std_logic;
    rematch009_in_chars              : in  std_logic_vector(31 downto 0);
    rematch009_in_chars_count        : in  std_logic_vector(2 downto 0);
    rematch009_in_unl_valid          : in  std_logic;
    rematch009_in_unl_ready          : out std_logic;
    rematch009_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch009_in_cmd_valid          : out std_logic;
    rematch009_in_cmd_ready          : in  std_logic;
    rematch009_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch009_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch009_in_cmd_ctrl           : out std_logic_vector(REMATCH009_IN_BUS_ADDR_WIDTH*2-1 downto 0);
    rematch009_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch010_in_valid              : in  std_logic;
    rematch010_in_ready              : out std_logic;
    rematch010_in_dvalid             : in  std_logic;
    rematch010_in_last               : in  std_logic;
    rematch010_in_length             : in  std_logic_vector(31 downto 0);
    rematch010_in_count              : in  std_logic_vector(0 downto 0);
    rematch010_in_chars_valid        : in  std_logic;
    rematch010_in_chars_ready        : out std_logic;
    rematch010_in_chars_dvalid       : in  std_logic;
    rematch010_in_chars_last         : in  std_logic;
    rematch010_in_chars              : in  std_logic_vector(31 downto 0);
    rematch010_in_chars_count        : in  std_logic_vector(2 downto 0);
    rematch010_in_unl_valid          : in  std_logic;
    rematch010_in_unl_ready          : out std_logic;
    rematch010_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch010_in_cmd_valid          : out std_logic;
    rematch010_in_cmd_ready          : in  std_logic;
    rematch010_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch010_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch010_in_cmd_ctrl           : out std_logic_vector(REMATCH010_IN_BUS_ADDR_WIDTH*2-1 downto 0);
    rematch010_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch011_in_valid              : in  std_logic;
    rematch011_in_ready              : out std_logic;
    rematch011_in_dvalid             : in  std_logic;
    rematch011_in_last               : in  std_logic;
    rematch011_in_length             : in  std_logic_vector(31 downto 0);
    rematch011_in_count              : in  std_logic_vector(0 downto 0);
    rematch011_in_chars_valid        : in  std_logic;
    rematch011_in_chars_ready        : out std_logic;
    rematch011_in_chars_dvalid       : in  std_logic;
    rematch011_in_chars_last         : in  std_logic;
    rematch011_in_chars              : in  std_logic_vector(31 downto 0);
    rematch011_in_chars_count        : in  std_logic_vector(2 downto 0);
    rematch011_in_unl_valid          : in  std_logic;
    rematch011_in_unl_ready          : out std_logic;
    rematch011_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch011_in_cmd_valid          : out std_logic;
    rematch011_in_cmd_ready          : in  std_logic;
    rematch011_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch011_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch011_in_cmd_ctrl           : out std_logic_vector(REMATCH011_IN_BUS_ADDR_WIDTH*2-1 downto 0);
    rematch011_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch012_in_valid              : in  std_logic;
    rematch012_in_ready              : out std_logic;
    rematch012_in_dvalid             : in  std_logic;
    rematch012_in_last               : in  std_logic;
    rematch012_in_length             : in  std_logic_vector(31 downto 0);
    rematch012_in_count              : in  std_logic_vector(0 downto 0);
    rematch012_in_chars_valid        : in  std_logic;
    rematch012_in_chars_ready        : out std_logic;
    rematch012_in_chars_dvalid       : in  std_logic;
    rematch012_in_chars_last         : in  std_logic;
    rematch012_in_chars              : in  std_logic_vector(31 downto 0);
    rematch012_in_chars_count        : in  std_logic_vector(2 downto 0);
    rematch012_in_unl_valid          : in  std_logic;
    rematch012_in_unl_ready          : out std_logic;
    rematch012_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch012_in_cmd_valid          : out std_logic;
    rematch012_in_cmd_ready          : in  std_logic;
    rematch012_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch012_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch012_in_cmd_ctrl           : out std_logic_vector(REMATCH012_IN_BUS_ADDR_WIDTH*2-1 downto 0);
    rematch012_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch013_in_valid              : in  std_logic;
    rematch013_in_ready              : out std_logic;
    rematch013_in_dvalid             : in  std_logic;
    rematch013_in_last               : in  std_logic;
    rematch013_in_length             : in  std_logic_vector(31 downto 0);
    rematch013_in_count              : in  std_logic_vector(0 downto 0);
    rematch013_in_chars_valid        : in  std_logic;
    rematch013_in_chars_ready        : out std_logic;
    rematch013_in_chars_dvalid       : in  std_logic;
    rematch013_in_chars_last         : in  std_logic;
    rematch013_in_chars              : in  std_logic_vector(31 downto 0);
    rematch013_in_chars_count        : in  std_logic_vector(2 downto 0);
    rematch013_in_unl_valid          : in  std_logic;
    rematch013_in_unl_ready          : out std_logic;
    rematch013_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch013_in_cmd_valid          : out std_logic;
    rematch013_in_cmd_ready          : in  std_logic;
    rematch013_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch013_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch013_in_cmd_ctrl           : out std_logic_vector(REMATCH013_IN_BUS_ADDR_WIDTH*2-1 downto 0);
    rematch013_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch014_in_valid              : in  std_logic;
    rematch014_in_ready              : out std_logic;
    rematch014_in_dvalid             : in  std_logic;
    rematch014_in_last               : in  std_logic;
    rematch014_in_length             : in  std_logic_vector(31 downto 0);
    rematch014_in_count              : in  std_logic_vector(0 downto 0);
    rematch014_in_chars_valid        : in  std_logic;
    rematch014_in_chars_ready        : out std_logic;
    rematch014_in_chars_dvalid       : in  std_logic;
    rematch014_in_chars_last         : in  std_logic;
    rematch014_in_chars              : in  std_logic_vector(31 downto 0);
    rematch014_in_chars_count        : in  std_logic_vector(2 downto 0);
    rematch014_in_unl_valid          : in  std_logic;
    rematch014_in_unl_ready          : out std_logic;
    rematch014_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch014_in_cmd_valid          : out std_logic;
    rematch014_in_cmd_ready          : in  std_logic;
    rematch014_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch014_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch014_in_cmd_ctrl           : out std_logic_vector(REMATCH014_IN_BUS_ADDR_WIDTH*2-1 downto 0);
    rematch014_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch015_in_valid              : in  std_logic;
    rematch015_in_ready              : out std_logic;
    rematch015_in_dvalid             : in  std_logic;
    rematch015_in_last               : in  std_logic;
    rematch015_in_length             : in  std_logic_vector(31 downto 0);
    rematch015_in_count              : in  std_logic_vector(0 downto 0);
    rematch015_in_chars_valid        : in  std_logic;
    rematch015_in_chars_ready        : out std_logic;
    rematch015_in_chars_dvalid       : in  std_logic;
    rematch015_in_chars_last         : in  std_logic;
    rematch015_in_chars              : in  std_logic_vector(31 downto 0);
    rematch015_in_chars_count        : in  std_logic_vector(2 downto 0);
    rematch015_in_unl_valid          : in  std_logic;
    rematch015_in_unl_ready          : out std_logic;
    rematch015_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch015_in_cmd_valid          : out std_logic;
    rematch015_in_cmd_ready          : in  std_logic;
    rematch015_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch015_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch015_in_cmd_ctrl           : out std_logic_vector(REMATCH015_IN_BUS_ADDR_WIDTH*2-1 downto 0);
    rematch015_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch000_taxi_out_valid        : out std_logic;
    rematch000_taxi_out_ready        : in  std_logic;
    rematch000_taxi_out_dvalid       : out std_logic;
    rematch000_taxi_out_last         : out std_logic;
    rematch000_taxi_out              : out std_logic_vector(31 downto 0);
    rematch000_taxi_out_unl_valid    : in  std_logic;
    rematch000_taxi_out_unl_ready    : out std_logic;
    rematch000_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch000_taxi_out_cmd_valid    : out std_logic;
    rematch000_taxi_out_cmd_ready    : in  std_logic;
    rematch000_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch000_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch000_taxi_out_cmd_ctrl     : out std_logic_vector(REMATCH000_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
    rematch000_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch001_taxi_out_valid        : out std_logic;
    rematch001_taxi_out_ready        : in  std_logic;
    rematch001_taxi_out_dvalid       : out std_logic;
    rematch001_taxi_out_last         : out std_logic;
    rematch001_taxi_out              : out std_logic_vector(31 downto 0);
    rematch001_taxi_out_unl_valid    : in  std_logic;
    rematch001_taxi_out_unl_ready    : out std_logic;
    rematch001_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch001_taxi_out_cmd_valid    : out std_logic;
    rematch001_taxi_out_cmd_ready    : in  std_logic;
    rematch001_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch001_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch001_taxi_out_cmd_ctrl     : out std_logic_vector(REMATCH001_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
    rematch001_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch002_taxi_out_valid        : out std_logic;
    rematch002_taxi_out_ready        : in  std_logic;
    rematch002_taxi_out_dvalid       : out std_logic;
    rematch002_taxi_out_last         : out std_logic;
    rematch002_taxi_out              : out std_logic_vector(31 downto 0);
    rematch002_taxi_out_unl_valid    : in  std_logic;
    rematch002_taxi_out_unl_ready    : out std_logic;
    rematch002_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch002_taxi_out_cmd_valid    : out std_logic;
    rematch002_taxi_out_cmd_ready    : in  std_logic;
    rematch002_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch002_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch002_taxi_out_cmd_ctrl     : out std_logic_vector(REMATCH002_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
    rematch002_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch003_taxi_out_valid        : out std_logic;
    rematch003_taxi_out_ready        : in  std_logic;
    rematch003_taxi_out_dvalid       : out std_logic;
    rematch003_taxi_out_last         : out std_logic;
    rematch003_taxi_out              : out std_logic_vector(31 downto 0);
    rematch003_taxi_out_unl_valid    : in  std_logic;
    rematch003_taxi_out_unl_ready    : out std_logic;
    rematch003_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch003_taxi_out_cmd_valid    : out std_logic;
    rematch003_taxi_out_cmd_ready    : in  std_logic;
    rematch003_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch003_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch003_taxi_out_cmd_ctrl     : out std_logic_vector(REMATCH003_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
    rematch003_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch004_taxi_out_valid        : out std_logic;
    rematch004_taxi_out_ready        : in  std_logic;
    rematch004_taxi_out_dvalid       : out std_logic;
    rematch004_taxi_out_last         : out std_logic;
    rematch004_taxi_out              : out std_logic_vector(31 downto 0);
    rematch004_taxi_out_unl_valid    : in  std_logic;
    rematch004_taxi_out_unl_ready    : out std_logic;
    rematch004_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch004_taxi_out_cmd_valid    : out std_logic;
    rematch004_taxi_out_cmd_ready    : in  std_logic;
    rematch004_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch004_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch004_taxi_out_cmd_ctrl     : out std_logic_vector(REMATCH004_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
    rematch004_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch005_taxi_out_valid        : out std_logic;
    rematch005_taxi_out_ready        : in  std_logic;
    rematch005_taxi_out_dvalid       : out std_logic;
    rematch005_taxi_out_last         : out std_logic;
    rematch005_taxi_out              : out std_logic_vector(31 downto 0);
    rematch005_taxi_out_unl_valid    : in  std_logic;
    rematch005_taxi_out_unl_ready    : out std_logic;
    rematch005_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch005_taxi_out_cmd_valid    : out std_logic;
    rematch005_taxi_out_cmd_ready    : in  std_logic;
    rematch005_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch005_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch005_taxi_out_cmd_ctrl     : out std_logic_vector(REMATCH005_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
    rematch005_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch006_taxi_out_valid        : out std_logic;
    rematch006_taxi_out_ready        : in  std_logic;
    rematch006_taxi_out_dvalid       : out std_logic;
    rematch006_taxi_out_last         : out std_logic;
    rematch006_taxi_out              : out std_logic_vector(31 downto 0);
    rematch006_taxi_out_unl_valid    : in  std_logic;
    rematch006_taxi_out_unl_ready    : out std_logic;
    rematch006_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch006_taxi_out_cmd_valid    : out std_logic;
    rematch006_taxi_out_cmd_ready    : in  std_logic;
    rematch006_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch006_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch006_taxi_out_cmd_ctrl     : out std_logic_vector(REMATCH006_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
    rematch006_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch007_taxi_out_valid        : out std_logic;
    rematch007_taxi_out_ready        : in  std_logic;
    rematch007_taxi_out_dvalid       : out std_logic;
    rematch007_taxi_out_last         : out std_logic;
    rematch007_taxi_out              : out std_logic_vector(31 downto 0);
    rematch007_taxi_out_unl_valid    : in  std_logic;
    rematch007_taxi_out_unl_ready    : out std_logic;
    rematch007_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch007_taxi_out_cmd_valid    : out std_logic;
    rematch007_taxi_out_cmd_ready    : in  std_logic;
    rematch007_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch007_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch007_taxi_out_cmd_ctrl     : out std_logic_vector(REMATCH007_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
    rematch007_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch008_taxi_out_valid        : out std_logic;
    rematch008_taxi_out_ready        : in  std_logic;
    rematch008_taxi_out_dvalid       : out std_logic;
    rematch008_taxi_out_last         : out std_logic;
    rematch008_taxi_out              : out std_logic_vector(31 downto 0);
    rematch008_taxi_out_unl_valid    : in  std_logic;
    rematch008_taxi_out_unl_ready    : out std_logic;
    rematch008_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch008_taxi_out_cmd_valid    : out std_logic;
    rematch008_taxi_out_cmd_ready    : in  std_logic;
    rematch008_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch008_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch008_taxi_out_cmd_ctrl     : out std_logic_vector(REMATCH008_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
    rematch008_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch009_taxi_out_valid        : out std_logic;
    rematch009_taxi_out_ready        : in  std_logic;
    rematch009_taxi_out_dvalid       : out std_logic;
    rematch009_taxi_out_last         : out std_logic;
    rematch009_taxi_out              : out std_logic_vector(31 downto 0);
    rematch009_taxi_out_unl_valid    : in  std_logic;
    rematch009_taxi_out_unl_ready    : out std_logic;
    rematch009_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch009_taxi_out_cmd_valid    : out std_logic;
    rematch009_taxi_out_cmd_ready    : in  std_logic;
    rematch009_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch009_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch009_taxi_out_cmd_ctrl     : out std_logic_vector(REMATCH009_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
    rematch009_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch010_taxi_out_valid        : out std_logic;
    rematch010_taxi_out_ready        : in  std_logic;
    rematch010_taxi_out_dvalid       : out std_logic;
    rematch010_taxi_out_last         : out std_logic;
    rematch010_taxi_out              : out std_logic_vector(31 downto 0);
    rematch010_taxi_out_unl_valid    : in  std_logic;
    rematch010_taxi_out_unl_ready    : out std_logic;
    rematch010_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch010_taxi_out_cmd_valid    : out std_logic;
    rematch010_taxi_out_cmd_ready    : in  std_logic;
    rematch010_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch010_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch010_taxi_out_cmd_ctrl     : out std_logic_vector(REMATCH010_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
    rematch010_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch011_taxi_out_valid        : out std_logic;
    rematch011_taxi_out_ready        : in  std_logic;
    rematch011_taxi_out_dvalid       : out std_logic;
    rematch011_taxi_out_last         : out std_logic;
    rematch011_taxi_out              : out std_logic_vector(31 downto 0);
    rematch011_taxi_out_unl_valid    : in  std_logic;
    rematch011_taxi_out_unl_ready    : out std_logic;
    rematch011_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch011_taxi_out_cmd_valid    : out std_logic;
    rematch011_taxi_out_cmd_ready    : in  std_logic;
    rematch011_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch011_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch011_taxi_out_cmd_ctrl     : out std_logic_vector(REMATCH011_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
    rematch011_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch012_taxi_out_valid        : out std_logic;
    rematch012_taxi_out_ready        : in  std_logic;
    rematch012_taxi_out_dvalid       : out std_logic;
    rematch012_taxi_out_last         : out std_logic;
    rematch012_taxi_out              : out std_logic_vector(31 downto 0);
    rematch012_taxi_out_unl_valid    : in  std_logic;
    rematch012_taxi_out_unl_ready    : out std_logic;
    rematch012_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch012_taxi_out_cmd_valid    : out std_logic;
    rematch012_taxi_out_cmd_ready    : in  std_logic;
    rematch012_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch012_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch012_taxi_out_cmd_ctrl     : out std_logic_vector(REMATCH012_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
    rematch012_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch013_taxi_out_valid        : out std_logic;
    rematch013_taxi_out_ready        : in  std_logic;
    rematch013_taxi_out_dvalid       : out std_logic;
    rematch013_taxi_out_last         : out std_logic;
    rematch013_taxi_out              : out std_logic_vector(31 downto 0);
    rematch013_taxi_out_unl_valid    : in  std_logic;
    rematch013_taxi_out_unl_ready    : out std_logic;
    rematch013_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch013_taxi_out_cmd_valid    : out std_logic;
    rematch013_taxi_out_cmd_ready    : in  std_logic;
    rematch013_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch013_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch013_taxi_out_cmd_ctrl     : out std_logic_vector(REMATCH013_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
    rematch013_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch014_taxi_out_valid        : out std_logic;
    rematch014_taxi_out_ready        : in  std_logic;
    rematch014_taxi_out_dvalid       : out std_logic;
    rematch014_taxi_out_last         : out std_logic;
    rematch014_taxi_out              : out std_logic_vector(31 downto 0);
    rematch014_taxi_out_unl_valid    : in  std_logic;
    rematch014_taxi_out_unl_ready    : out std_logic;
    rematch014_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch014_taxi_out_cmd_valid    : out std_logic;
    rematch014_taxi_out_cmd_ready    : in  std_logic;
    rematch014_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch014_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch014_taxi_out_cmd_ctrl     : out std_logic_vector(REMATCH014_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
    rematch014_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch015_taxi_out_valid        : out std_logic;
    rematch015_taxi_out_ready        : in  std_logic;
    rematch015_taxi_out_dvalid       : out std_logic;
    rematch015_taxi_out_last         : out std_logic;
    rematch015_taxi_out              : out std_logic_vector(31 downto 0);
    rematch015_taxi_out_unl_valid    : in  std_logic;
    rematch015_taxi_out_unl_ready    : out std_logic;
    rematch015_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    rematch015_taxi_out_cmd_valid    : out std_logic;
    rematch015_taxi_out_cmd_ready    : in  std_logic;
    rematch015_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch015_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    rematch015_taxi_out_cmd_ctrl     : out std_logic_vector(REMATCH015_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
    rematch015_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0)
  );
end entity;

architecture Implementation of Kernel_Nucleus is
  component Kernel is
    generic (
      INDEX_WIDTH : integer := 32;
      TAG_WIDTH   : integer := 1
    );
    port (
      kcd_clk                          : in  std_logic;
      kcd_reset                        : in  std_logic;
      rematch000_in_valid              : in  std_logic;
      rematch000_in_ready              : out std_logic;
      rematch000_in_dvalid             : in  std_logic;
      rematch000_in_last               : in  std_logic;
      rematch000_in_length             : in  std_logic_vector(31 downto 0);
      rematch000_in_count              : in  std_logic_vector(0 downto 0);
      rematch000_in_chars_valid        : in  std_logic;
      rematch000_in_chars_ready        : out std_logic;
      rematch000_in_chars_dvalid       : in  std_logic;
      rematch000_in_chars_last         : in  std_logic;
      rematch000_in_chars              : in  std_logic_vector(31 downto 0);
      rematch000_in_chars_count        : in  std_logic_vector(2 downto 0);
      rematch000_in_unl_valid          : in  std_logic;
      rematch000_in_unl_ready          : out std_logic;
      rematch000_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch000_in_cmd_valid          : out std_logic;
      rematch000_in_cmd_ready          : in  std_logic;
      rematch000_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch000_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch000_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch001_in_valid              : in  std_logic;
      rematch001_in_ready              : out std_logic;
      rematch001_in_dvalid             : in  std_logic;
      rematch001_in_last               : in  std_logic;
      rematch001_in_length             : in  std_logic_vector(31 downto 0);
      rematch001_in_count              : in  std_logic_vector(0 downto 0);
      rematch001_in_chars_valid        : in  std_logic;
      rematch001_in_chars_ready        : out std_logic;
      rematch001_in_chars_dvalid       : in  std_logic;
      rematch001_in_chars_last         : in  std_logic;
      rematch001_in_chars              : in  std_logic_vector(31 downto 0);
      rematch001_in_chars_count        : in  std_logic_vector(2 downto 0);
      rematch001_in_unl_valid          : in  std_logic;
      rematch001_in_unl_ready          : out std_logic;
      rematch001_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch001_in_cmd_valid          : out std_logic;
      rematch001_in_cmd_ready          : in  std_logic;
      rematch001_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch001_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch001_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch002_in_valid              : in  std_logic;
      rematch002_in_ready              : out std_logic;
      rematch002_in_dvalid             : in  std_logic;
      rematch002_in_last               : in  std_logic;
      rematch002_in_length             : in  std_logic_vector(31 downto 0);
      rematch002_in_count              : in  std_logic_vector(0 downto 0);
      rematch002_in_chars_valid        : in  std_logic;
      rematch002_in_chars_ready        : out std_logic;
      rematch002_in_chars_dvalid       : in  std_logic;
      rematch002_in_chars_last         : in  std_logic;
      rematch002_in_chars              : in  std_logic_vector(31 downto 0);
      rematch002_in_chars_count        : in  std_logic_vector(2 downto 0);
      rematch002_in_unl_valid          : in  std_logic;
      rematch002_in_unl_ready          : out std_logic;
      rematch002_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch002_in_cmd_valid          : out std_logic;
      rematch002_in_cmd_ready          : in  std_logic;
      rematch002_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch002_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch002_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch003_in_valid              : in  std_logic;
      rematch003_in_ready              : out std_logic;
      rematch003_in_dvalid             : in  std_logic;
      rematch003_in_last               : in  std_logic;
      rematch003_in_length             : in  std_logic_vector(31 downto 0);
      rematch003_in_count              : in  std_logic_vector(0 downto 0);
      rematch003_in_chars_valid        : in  std_logic;
      rematch003_in_chars_ready        : out std_logic;
      rematch003_in_chars_dvalid       : in  std_logic;
      rematch003_in_chars_last         : in  std_logic;
      rematch003_in_chars              : in  std_logic_vector(31 downto 0);
      rematch003_in_chars_count        : in  std_logic_vector(2 downto 0);
      rematch003_in_unl_valid          : in  std_logic;
      rematch003_in_unl_ready          : out std_logic;
      rematch003_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch003_in_cmd_valid          : out std_logic;
      rematch003_in_cmd_ready          : in  std_logic;
      rematch003_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch003_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch003_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch004_in_valid              : in  std_logic;
      rematch004_in_ready              : out std_logic;
      rematch004_in_dvalid             : in  std_logic;
      rematch004_in_last               : in  std_logic;
      rematch004_in_length             : in  std_logic_vector(31 downto 0);
      rematch004_in_count              : in  std_logic_vector(0 downto 0);
      rematch004_in_chars_valid        : in  std_logic;
      rematch004_in_chars_ready        : out std_logic;
      rematch004_in_chars_dvalid       : in  std_logic;
      rematch004_in_chars_last         : in  std_logic;
      rematch004_in_chars              : in  std_logic_vector(31 downto 0);
      rematch004_in_chars_count        : in  std_logic_vector(2 downto 0);
      rematch004_in_unl_valid          : in  std_logic;
      rematch004_in_unl_ready          : out std_logic;
      rematch004_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch004_in_cmd_valid          : out std_logic;
      rematch004_in_cmd_ready          : in  std_logic;
      rematch004_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch004_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch004_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch005_in_valid              : in  std_logic;
      rematch005_in_ready              : out std_logic;
      rematch005_in_dvalid             : in  std_logic;
      rematch005_in_last               : in  std_logic;
      rematch005_in_length             : in  std_logic_vector(31 downto 0);
      rematch005_in_count              : in  std_logic_vector(0 downto 0);
      rematch005_in_chars_valid        : in  std_logic;
      rematch005_in_chars_ready        : out std_logic;
      rematch005_in_chars_dvalid       : in  std_logic;
      rematch005_in_chars_last         : in  std_logic;
      rematch005_in_chars              : in  std_logic_vector(31 downto 0);
      rematch005_in_chars_count        : in  std_logic_vector(2 downto 0);
      rematch005_in_unl_valid          : in  std_logic;
      rematch005_in_unl_ready          : out std_logic;
      rematch005_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch005_in_cmd_valid          : out std_logic;
      rematch005_in_cmd_ready          : in  std_logic;
      rematch005_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch005_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch005_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch006_in_valid              : in  std_logic;
      rematch006_in_ready              : out std_logic;
      rematch006_in_dvalid             : in  std_logic;
      rematch006_in_last               : in  std_logic;
      rematch006_in_length             : in  std_logic_vector(31 downto 0);
      rematch006_in_count              : in  std_logic_vector(0 downto 0);
      rematch006_in_chars_valid        : in  std_logic;
      rematch006_in_chars_ready        : out std_logic;
      rematch006_in_chars_dvalid       : in  std_logic;
      rematch006_in_chars_last         : in  std_logic;
      rematch006_in_chars              : in  std_logic_vector(31 downto 0);
      rematch006_in_chars_count        : in  std_logic_vector(2 downto 0);
      rematch006_in_unl_valid          : in  std_logic;
      rematch006_in_unl_ready          : out std_logic;
      rematch006_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch006_in_cmd_valid          : out std_logic;
      rematch006_in_cmd_ready          : in  std_logic;
      rematch006_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch006_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch006_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch007_in_valid              : in  std_logic;
      rematch007_in_ready              : out std_logic;
      rematch007_in_dvalid             : in  std_logic;
      rematch007_in_last               : in  std_logic;
      rematch007_in_length             : in  std_logic_vector(31 downto 0);
      rematch007_in_count              : in  std_logic_vector(0 downto 0);
      rematch007_in_chars_valid        : in  std_logic;
      rematch007_in_chars_ready        : out std_logic;
      rematch007_in_chars_dvalid       : in  std_logic;
      rematch007_in_chars_last         : in  std_logic;
      rematch007_in_chars              : in  std_logic_vector(31 downto 0);
      rematch007_in_chars_count        : in  std_logic_vector(2 downto 0);
      rematch007_in_unl_valid          : in  std_logic;
      rematch007_in_unl_ready          : out std_logic;
      rematch007_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch007_in_cmd_valid          : out std_logic;
      rematch007_in_cmd_ready          : in  std_logic;
      rematch007_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch007_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch007_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch008_in_valid              : in  std_logic;
      rematch008_in_ready              : out std_logic;
      rematch008_in_dvalid             : in  std_logic;
      rematch008_in_last               : in  std_logic;
      rematch008_in_length             : in  std_logic_vector(31 downto 0);
      rematch008_in_count              : in  std_logic_vector(0 downto 0);
      rematch008_in_chars_valid        : in  std_logic;
      rematch008_in_chars_ready        : out std_logic;
      rematch008_in_chars_dvalid       : in  std_logic;
      rematch008_in_chars_last         : in  std_logic;
      rematch008_in_chars              : in  std_logic_vector(31 downto 0);
      rematch008_in_chars_count        : in  std_logic_vector(2 downto 0);
      rematch008_in_unl_valid          : in  std_logic;
      rematch008_in_unl_ready          : out std_logic;
      rematch008_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch008_in_cmd_valid          : out std_logic;
      rematch008_in_cmd_ready          : in  std_logic;
      rematch008_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch008_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch008_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch009_in_valid              : in  std_logic;
      rematch009_in_ready              : out std_logic;
      rematch009_in_dvalid             : in  std_logic;
      rematch009_in_last               : in  std_logic;
      rematch009_in_length             : in  std_logic_vector(31 downto 0);
      rematch009_in_count              : in  std_logic_vector(0 downto 0);
      rematch009_in_chars_valid        : in  std_logic;
      rematch009_in_chars_ready        : out std_logic;
      rematch009_in_chars_dvalid       : in  std_logic;
      rematch009_in_chars_last         : in  std_logic;
      rematch009_in_chars              : in  std_logic_vector(31 downto 0);
      rematch009_in_chars_count        : in  std_logic_vector(2 downto 0);
      rematch009_in_unl_valid          : in  std_logic;
      rematch009_in_unl_ready          : out std_logic;
      rematch009_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch009_in_cmd_valid          : out std_logic;
      rematch009_in_cmd_ready          : in  std_logic;
      rematch009_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch009_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch009_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch010_in_valid              : in  std_logic;
      rematch010_in_ready              : out std_logic;
      rematch010_in_dvalid             : in  std_logic;
      rematch010_in_last               : in  std_logic;
      rematch010_in_length             : in  std_logic_vector(31 downto 0);
      rematch010_in_count              : in  std_logic_vector(0 downto 0);
      rematch010_in_chars_valid        : in  std_logic;
      rematch010_in_chars_ready        : out std_logic;
      rematch010_in_chars_dvalid       : in  std_logic;
      rematch010_in_chars_last         : in  std_logic;
      rematch010_in_chars              : in  std_logic_vector(31 downto 0);
      rematch010_in_chars_count        : in  std_logic_vector(2 downto 0);
      rematch010_in_unl_valid          : in  std_logic;
      rematch010_in_unl_ready          : out std_logic;
      rematch010_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch010_in_cmd_valid          : out std_logic;
      rematch010_in_cmd_ready          : in  std_logic;
      rematch010_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch010_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch010_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch011_in_valid              : in  std_logic;
      rematch011_in_ready              : out std_logic;
      rematch011_in_dvalid             : in  std_logic;
      rematch011_in_last               : in  std_logic;
      rematch011_in_length             : in  std_logic_vector(31 downto 0);
      rematch011_in_count              : in  std_logic_vector(0 downto 0);
      rematch011_in_chars_valid        : in  std_logic;
      rematch011_in_chars_ready        : out std_logic;
      rematch011_in_chars_dvalid       : in  std_logic;
      rematch011_in_chars_last         : in  std_logic;
      rematch011_in_chars              : in  std_logic_vector(31 downto 0);
      rematch011_in_chars_count        : in  std_logic_vector(2 downto 0);
      rematch011_in_unl_valid          : in  std_logic;
      rematch011_in_unl_ready          : out std_logic;
      rematch011_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch011_in_cmd_valid          : out std_logic;
      rematch011_in_cmd_ready          : in  std_logic;
      rematch011_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch011_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch011_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch012_in_valid              : in  std_logic;
      rematch012_in_ready              : out std_logic;
      rematch012_in_dvalid             : in  std_logic;
      rematch012_in_last               : in  std_logic;
      rematch012_in_length             : in  std_logic_vector(31 downto 0);
      rematch012_in_count              : in  std_logic_vector(0 downto 0);
      rematch012_in_chars_valid        : in  std_logic;
      rematch012_in_chars_ready        : out std_logic;
      rematch012_in_chars_dvalid       : in  std_logic;
      rematch012_in_chars_last         : in  std_logic;
      rematch012_in_chars              : in  std_logic_vector(31 downto 0);
      rematch012_in_chars_count        : in  std_logic_vector(2 downto 0);
      rematch012_in_unl_valid          : in  std_logic;
      rematch012_in_unl_ready          : out std_logic;
      rematch012_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch012_in_cmd_valid          : out std_logic;
      rematch012_in_cmd_ready          : in  std_logic;
      rematch012_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch012_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch012_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch013_in_valid              : in  std_logic;
      rematch013_in_ready              : out std_logic;
      rematch013_in_dvalid             : in  std_logic;
      rematch013_in_last               : in  std_logic;
      rematch013_in_length             : in  std_logic_vector(31 downto 0);
      rematch013_in_count              : in  std_logic_vector(0 downto 0);
      rematch013_in_chars_valid        : in  std_logic;
      rematch013_in_chars_ready        : out std_logic;
      rematch013_in_chars_dvalid       : in  std_logic;
      rematch013_in_chars_last         : in  std_logic;
      rematch013_in_chars              : in  std_logic_vector(31 downto 0);
      rematch013_in_chars_count        : in  std_logic_vector(2 downto 0);
      rematch013_in_unl_valid          : in  std_logic;
      rematch013_in_unl_ready          : out std_logic;
      rematch013_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch013_in_cmd_valid          : out std_logic;
      rematch013_in_cmd_ready          : in  std_logic;
      rematch013_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch013_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch013_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch014_in_valid              : in  std_logic;
      rematch014_in_ready              : out std_logic;
      rematch014_in_dvalid             : in  std_logic;
      rematch014_in_last               : in  std_logic;
      rematch014_in_length             : in  std_logic_vector(31 downto 0);
      rematch014_in_count              : in  std_logic_vector(0 downto 0);
      rematch014_in_chars_valid        : in  std_logic;
      rematch014_in_chars_ready        : out std_logic;
      rematch014_in_chars_dvalid       : in  std_logic;
      rematch014_in_chars_last         : in  std_logic;
      rematch014_in_chars              : in  std_logic_vector(31 downto 0);
      rematch014_in_chars_count        : in  std_logic_vector(2 downto 0);
      rematch014_in_unl_valid          : in  std_logic;
      rematch014_in_unl_ready          : out std_logic;
      rematch014_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch014_in_cmd_valid          : out std_logic;
      rematch014_in_cmd_ready          : in  std_logic;
      rematch014_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch014_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch014_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch015_in_valid              : in  std_logic;
      rematch015_in_ready              : out std_logic;
      rematch015_in_dvalid             : in  std_logic;
      rematch015_in_last               : in  std_logic;
      rematch015_in_length             : in  std_logic_vector(31 downto 0);
      rematch015_in_count              : in  std_logic_vector(0 downto 0);
      rematch015_in_chars_valid        : in  std_logic;
      rematch015_in_chars_ready        : out std_logic;
      rematch015_in_chars_dvalid       : in  std_logic;
      rematch015_in_chars_last         : in  std_logic;
      rematch015_in_chars              : in  std_logic_vector(31 downto 0);
      rematch015_in_chars_count        : in  std_logic_vector(2 downto 0);
      rematch015_in_unl_valid          : in  std_logic;
      rematch015_in_unl_ready          : out std_logic;
      rematch015_in_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch015_in_cmd_valid          : out std_logic;
      rematch015_in_cmd_ready          : in  std_logic;
      rematch015_in_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch015_in_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch015_in_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch000_taxi_out_valid        : out std_logic;
      rematch000_taxi_out_ready        : in  std_logic;
      rematch000_taxi_out_dvalid       : out std_logic;
      rematch000_taxi_out_last         : out std_logic;
      rematch000_taxi_out              : out std_logic_vector(31 downto 0);
      rematch000_taxi_out_unl_valid    : in  std_logic;
      rematch000_taxi_out_unl_ready    : out std_logic;
      rematch000_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch000_taxi_out_cmd_valid    : out std_logic;
      rematch000_taxi_out_cmd_ready    : in  std_logic;
      rematch000_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch000_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch000_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch001_taxi_out_valid        : out std_logic;
      rematch001_taxi_out_ready        : in  std_logic;
      rematch001_taxi_out_dvalid       : out std_logic;
      rematch001_taxi_out_last         : out std_logic;
      rematch001_taxi_out              : out std_logic_vector(31 downto 0);
      rematch001_taxi_out_unl_valid    : in  std_logic;
      rematch001_taxi_out_unl_ready    : out std_logic;
      rematch001_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch001_taxi_out_cmd_valid    : out std_logic;
      rematch001_taxi_out_cmd_ready    : in  std_logic;
      rematch001_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch001_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch001_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch002_taxi_out_valid        : out std_logic;
      rematch002_taxi_out_ready        : in  std_logic;
      rematch002_taxi_out_dvalid       : out std_logic;
      rematch002_taxi_out_last         : out std_logic;
      rematch002_taxi_out              : out std_logic_vector(31 downto 0);
      rematch002_taxi_out_unl_valid    : in  std_logic;
      rematch002_taxi_out_unl_ready    : out std_logic;
      rematch002_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch002_taxi_out_cmd_valid    : out std_logic;
      rematch002_taxi_out_cmd_ready    : in  std_logic;
      rematch002_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch002_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch002_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch003_taxi_out_valid        : out std_logic;
      rematch003_taxi_out_ready        : in  std_logic;
      rematch003_taxi_out_dvalid       : out std_logic;
      rematch003_taxi_out_last         : out std_logic;
      rematch003_taxi_out              : out std_logic_vector(31 downto 0);
      rematch003_taxi_out_unl_valid    : in  std_logic;
      rematch003_taxi_out_unl_ready    : out std_logic;
      rematch003_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch003_taxi_out_cmd_valid    : out std_logic;
      rematch003_taxi_out_cmd_ready    : in  std_logic;
      rematch003_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch003_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch003_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch004_taxi_out_valid        : out std_logic;
      rematch004_taxi_out_ready        : in  std_logic;
      rematch004_taxi_out_dvalid       : out std_logic;
      rematch004_taxi_out_last         : out std_logic;
      rematch004_taxi_out              : out std_logic_vector(31 downto 0);
      rematch004_taxi_out_unl_valid    : in  std_logic;
      rematch004_taxi_out_unl_ready    : out std_logic;
      rematch004_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch004_taxi_out_cmd_valid    : out std_logic;
      rematch004_taxi_out_cmd_ready    : in  std_logic;
      rematch004_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch004_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch004_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch005_taxi_out_valid        : out std_logic;
      rematch005_taxi_out_ready        : in  std_logic;
      rematch005_taxi_out_dvalid       : out std_logic;
      rematch005_taxi_out_last         : out std_logic;
      rematch005_taxi_out              : out std_logic_vector(31 downto 0);
      rematch005_taxi_out_unl_valid    : in  std_logic;
      rematch005_taxi_out_unl_ready    : out std_logic;
      rematch005_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch005_taxi_out_cmd_valid    : out std_logic;
      rematch005_taxi_out_cmd_ready    : in  std_logic;
      rematch005_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch005_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch005_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch006_taxi_out_valid        : out std_logic;
      rematch006_taxi_out_ready        : in  std_logic;
      rematch006_taxi_out_dvalid       : out std_logic;
      rematch006_taxi_out_last         : out std_logic;
      rematch006_taxi_out              : out std_logic_vector(31 downto 0);
      rematch006_taxi_out_unl_valid    : in  std_logic;
      rematch006_taxi_out_unl_ready    : out std_logic;
      rematch006_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch006_taxi_out_cmd_valid    : out std_logic;
      rematch006_taxi_out_cmd_ready    : in  std_logic;
      rematch006_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch006_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch006_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch007_taxi_out_valid        : out std_logic;
      rematch007_taxi_out_ready        : in  std_logic;
      rematch007_taxi_out_dvalid       : out std_logic;
      rematch007_taxi_out_last         : out std_logic;
      rematch007_taxi_out              : out std_logic_vector(31 downto 0);
      rematch007_taxi_out_unl_valid    : in  std_logic;
      rematch007_taxi_out_unl_ready    : out std_logic;
      rematch007_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch007_taxi_out_cmd_valid    : out std_logic;
      rematch007_taxi_out_cmd_ready    : in  std_logic;
      rematch007_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch007_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch007_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch008_taxi_out_valid        : out std_logic;
      rematch008_taxi_out_ready        : in  std_logic;
      rematch008_taxi_out_dvalid       : out std_logic;
      rematch008_taxi_out_last         : out std_logic;
      rematch008_taxi_out              : out std_logic_vector(31 downto 0);
      rematch008_taxi_out_unl_valid    : in  std_logic;
      rematch008_taxi_out_unl_ready    : out std_logic;
      rematch008_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch008_taxi_out_cmd_valid    : out std_logic;
      rematch008_taxi_out_cmd_ready    : in  std_logic;
      rematch008_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch008_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch008_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch009_taxi_out_valid        : out std_logic;
      rematch009_taxi_out_ready        : in  std_logic;
      rematch009_taxi_out_dvalid       : out std_logic;
      rematch009_taxi_out_last         : out std_logic;
      rematch009_taxi_out              : out std_logic_vector(31 downto 0);
      rematch009_taxi_out_unl_valid    : in  std_logic;
      rematch009_taxi_out_unl_ready    : out std_logic;
      rematch009_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch009_taxi_out_cmd_valid    : out std_logic;
      rematch009_taxi_out_cmd_ready    : in  std_logic;
      rematch009_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch009_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch009_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch010_taxi_out_valid        : out std_logic;
      rematch010_taxi_out_ready        : in  std_logic;
      rematch010_taxi_out_dvalid       : out std_logic;
      rematch010_taxi_out_last         : out std_logic;
      rematch010_taxi_out              : out std_logic_vector(31 downto 0);
      rematch010_taxi_out_unl_valid    : in  std_logic;
      rematch010_taxi_out_unl_ready    : out std_logic;
      rematch010_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch010_taxi_out_cmd_valid    : out std_logic;
      rematch010_taxi_out_cmd_ready    : in  std_logic;
      rematch010_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch010_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch010_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch011_taxi_out_valid        : out std_logic;
      rematch011_taxi_out_ready        : in  std_logic;
      rematch011_taxi_out_dvalid       : out std_logic;
      rematch011_taxi_out_last         : out std_logic;
      rematch011_taxi_out              : out std_logic_vector(31 downto 0);
      rematch011_taxi_out_unl_valid    : in  std_logic;
      rematch011_taxi_out_unl_ready    : out std_logic;
      rematch011_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch011_taxi_out_cmd_valid    : out std_logic;
      rematch011_taxi_out_cmd_ready    : in  std_logic;
      rematch011_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch011_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch011_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch012_taxi_out_valid        : out std_logic;
      rematch012_taxi_out_ready        : in  std_logic;
      rematch012_taxi_out_dvalid       : out std_logic;
      rematch012_taxi_out_last         : out std_logic;
      rematch012_taxi_out              : out std_logic_vector(31 downto 0);
      rematch012_taxi_out_unl_valid    : in  std_logic;
      rematch012_taxi_out_unl_ready    : out std_logic;
      rematch012_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch012_taxi_out_cmd_valid    : out std_logic;
      rematch012_taxi_out_cmd_ready    : in  std_logic;
      rematch012_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch012_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch012_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch013_taxi_out_valid        : out std_logic;
      rematch013_taxi_out_ready        : in  std_logic;
      rematch013_taxi_out_dvalid       : out std_logic;
      rematch013_taxi_out_last         : out std_logic;
      rematch013_taxi_out              : out std_logic_vector(31 downto 0);
      rematch013_taxi_out_unl_valid    : in  std_logic;
      rematch013_taxi_out_unl_ready    : out std_logic;
      rematch013_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch013_taxi_out_cmd_valid    : out std_logic;
      rematch013_taxi_out_cmd_ready    : in  std_logic;
      rematch013_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch013_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch013_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch014_taxi_out_valid        : out std_logic;
      rematch014_taxi_out_ready        : in  std_logic;
      rematch014_taxi_out_dvalid       : out std_logic;
      rematch014_taxi_out_last         : out std_logic;
      rematch014_taxi_out              : out std_logic_vector(31 downto 0);
      rematch014_taxi_out_unl_valid    : in  std_logic;
      rematch014_taxi_out_unl_ready    : out std_logic;
      rematch014_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch014_taxi_out_cmd_valid    : out std_logic;
      rematch014_taxi_out_cmd_ready    : in  std_logic;
      rematch014_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch014_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch014_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch015_taxi_out_valid        : out std_logic;
      rematch015_taxi_out_ready        : in  std_logic;
      rematch015_taxi_out_dvalid       : out std_logic;
      rematch015_taxi_out_last         : out std_logic;
      rematch015_taxi_out              : out std_logic_vector(31 downto 0);
      rematch015_taxi_out_unl_valid    : in  std_logic;
      rematch015_taxi_out_unl_ready    : out std_logic;
      rematch015_taxi_out_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch015_taxi_out_cmd_valid    : out std_logic;
      rematch015_taxi_out_cmd_ready    : in  std_logic;
      rematch015_taxi_out_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch015_taxi_out_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch015_taxi_out_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      start                            : in  std_logic;
      stop                             : in  std_logic;
      reset                            : in  std_logic;
      idle                             : out std_logic;
      busy                             : out std_logic;
      done                             : out std_logic;
      result                           : out std_logic_vector(63 downto 0);
      rematch000_firstidx              : in  std_logic_vector(31 downto 0);
      rematch000_lastidx               : in  std_logic_vector(31 downto 0);
      rematch001_firstidx              : in  std_logic_vector(31 downto 0);
      rematch001_lastidx               : in  std_logic_vector(31 downto 0);
      rematch002_firstidx              : in  std_logic_vector(31 downto 0);
      rematch002_lastidx               : in  std_logic_vector(31 downto 0);
      rematch003_firstidx              : in  std_logic_vector(31 downto 0);
      rematch003_lastidx               : in  std_logic_vector(31 downto 0);
      rematch004_firstidx              : in  std_logic_vector(31 downto 0);
      rematch004_lastidx               : in  std_logic_vector(31 downto 0);
      rematch005_firstidx              : in  std_logic_vector(31 downto 0);
      rematch005_lastidx               : in  std_logic_vector(31 downto 0);
      rematch006_firstidx              : in  std_logic_vector(31 downto 0);
      rematch006_lastidx               : in  std_logic_vector(31 downto 0);
      rematch007_firstidx              : in  std_logic_vector(31 downto 0);
      rematch007_lastidx               : in  std_logic_vector(31 downto 0);
      rematch008_firstidx              : in  std_logic_vector(31 downto 0);
      rematch008_lastidx               : in  std_logic_vector(31 downto 0);
      rematch009_firstidx              : in  std_logic_vector(31 downto 0);
      rematch009_lastidx               : in  std_logic_vector(31 downto 0);
      rematch010_firstidx              : in  std_logic_vector(31 downto 0);
      rematch010_lastidx               : in  std_logic_vector(31 downto 0);
      rematch011_firstidx              : in  std_logic_vector(31 downto 0);
      rematch011_lastidx               : in  std_logic_vector(31 downto 0);
      rematch012_firstidx              : in  std_logic_vector(31 downto 0);
      rematch012_lastidx               : in  std_logic_vector(31 downto 0);
      rematch013_firstidx              : in  std_logic_vector(31 downto 0);
      rematch013_lastidx               : in  std_logic_vector(31 downto 0);
      rematch014_firstidx              : in  std_logic_vector(31 downto 0);
      rematch014_lastidx               : in  std_logic_vector(31 downto 0);
      rematch015_firstidx              : in  std_logic_vector(31 downto 0);
      rematch015_lastidx               : in  std_logic_vector(31 downto 0);
      rematch000_taxi_firstidx         : in  std_logic_vector(31 downto 0);
      rematch000_taxi_lastidx          : in  std_logic_vector(31 downto 0);
      rematch001_taxi_firstidx         : in  std_logic_vector(31 downto 0);
      rematch001_taxi_lastidx          : in  std_logic_vector(31 downto 0);
      rematch002_taxi_firstidx         : in  std_logic_vector(31 downto 0);
      rematch002_taxi_lastidx          : in  std_logic_vector(31 downto 0);
      rematch003_taxi_firstidx         : in  std_logic_vector(31 downto 0);
      rematch003_taxi_lastidx          : in  std_logic_vector(31 downto 0);
      rematch004_taxi_firstidx         : in  std_logic_vector(31 downto 0);
      rematch004_taxi_lastidx          : in  std_logic_vector(31 downto 0);
      rematch005_taxi_firstidx         : in  std_logic_vector(31 downto 0);
      rematch005_taxi_lastidx          : in  std_logic_vector(31 downto 0);
      rematch006_taxi_firstidx         : in  std_logic_vector(31 downto 0);
      rematch006_taxi_lastidx          : in  std_logic_vector(31 downto 0);
      rematch007_taxi_firstidx         : in  std_logic_vector(31 downto 0);
      rematch007_taxi_lastidx          : in  std_logic_vector(31 downto 0);
      rematch008_taxi_firstidx         : in  std_logic_vector(31 downto 0);
      rematch008_taxi_lastidx          : in  std_logic_vector(31 downto 0);
      rematch009_taxi_firstidx         : in  std_logic_vector(31 downto 0);
      rematch009_taxi_lastidx          : in  std_logic_vector(31 downto 0);
      rematch010_taxi_firstidx         : in  std_logic_vector(31 downto 0);
      rematch010_taxi_lastidx          : in  std_logic_vector(31 downto 0);
      rematch011_taxi_firstidx         : in  std_logic_vector(31 downto 0);
      rematch011_taxi_lastidx          : in  std_logic_vector(31 downto 0);
      rematch012_taxi_firstidx         : in  std_logic_vector(31 downto 0);
      rematch012_taxi_lastidx          : in  std_logic_vector(31 downto 0);
      rematch013_taxi_firstidx         : in  std_logic_vector(31 downto 0);
      rematch013_taxi_lastidx          : in  std_logic_vector(31 downto 0);
      rematch014_taxi_firstidx         : in  std_logic_vector(31 downto 0);
      rematch014_taxi_lastidx          : in  std_logic_vector(31 downto 0);
      rematch015_taxi_firstidx         : in  std_logic_vector(31 downto 0);
      rematch015_taxi_lastidx          : in  std_logic_vector(31 downto 0);
      rematch000_taxi_count            : out std_logic_vector(31 downto 0);
      rematch000_errors                : out std_logic_vector(31 downto 0);
      rematch001_taxi_count            : out std_logic_vector(31 downto 0);
      rematch001_errors                : out std_logic_vector(31 downto 0);
      rematch002_taxi_count            : out std_logic_vector(31 downto 0);
      rematch002_errors                : out std_logic_vector(31 downto 0);
      rematch003_taxi_count            : out std_logic_vector(31 downto 0);
      rematch003_errors                : out std_logic_vector(31 downto 0);
      rematch004_taxi_count            : out std_logic_vector(31 downto 0);
      rematch004_errors                : out std_logic_vector(31 downto 0);
      rematch005_taxi_count            : out std_logic_vector(31 downto 0);
      rematch005_errors                : out std_logic_vector(31 downto 0);
      rematch006_taxi_count            : out std_logic_vector(31 downto 0);
      rematch006_errors                : out std_logic_vector(31 downto 0);
      rematch007_taxi_count            : out std_logic_vector(31 downto 0);
      rematch007_errors                : out std_logic_vector(31 downto 0);
      rematch008_taxi_count            : out std_logic_vector(31 downto 0);
      rematch008_errors                : out std_logic_vector(31 downto 0);
      rematch009_taxi_count            : out std_logic_vector(31 downto 0);
      rematch009_errors                : out std_logic_vector(31 downto 0);
      rematch010_taxi_count            : out std_logic_vector(31 downto 0);
      rematch010_errors                : out std_logic_vector(31 downto 0);
      rematch011_taxi_count            : out std_logic_vector(31 downto 0);
      rematch011_errors                : out std_logic_vector(31 downto 0);
      rematch012_taxi_count            : out std_logic_vector(31 downto 0);
      rematch012_errors                : out std_logic_vector(31 downto 0);
      rematch013_taxi_count            : out std_logic_vector(31 downto 0);
      rematch013_errors                : out std_logic_vector(31 downto 0);
      rematch014_taxi_count            : out std_logic_vector(31 downto 0);
      rematch014_errors                : out std_logic_vector(31 downto 0);
      rematch015_taxi_count            : out std_logic_vector(31 downto 0);
      rematch015_errors                : out std_logic_vector(31 downto 0)
    );
  end component;

  signal Kernel_inst_rematch000_in_valid                        : std_logic;
  signal Kernel_inst_rematch000_in_ready                        : std_logic;
  signal Kernel_inst_rematch000_in_dvalid                       : std_logic;
  signal Kernel_inst_rematch000_in_last                         : std_logic;
  signal Kernel_inst_rematch000_in_length                       : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch000_in_count                        : std_logic_vector(0 downto 0);
  signal Kernel_inst_rematch000_in_chars_valid                  : std_logic;
  signal Kernel_inst_rematch000_in_chars_ready                  : std_logic;
  signal Kernel_inst_rematch000_in_chars_dvalid                 : std_logic;
  signal Kernel_inst_rematch000_in_chars_last                   : std_logic;
  signal Kernel_inst_rematch000_in_chars                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch000_in_chars_count                  : std_logic_vector(2 downto 0);

  signal Kernel_inst_rematch000_in_unl_valid                    : std_logic;
  signal Kernel_inst_rematch000_in_unl_ready                    : std_logic;
  signal Kernel_inst_rematch000_in_unl_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch000_in_cmd_valid                    : std_logic;
  signal Kernel_inst_rematch000_in_cmd_ready                    : std_logic;
  signal Kernel_inst_rematch000_in_cmd_firstIdx                 : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch000_in_cmd_lastIdx                  : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch000_in_cmd_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch001_in_valid                        : std_logic;
  signal Kernel_inst_rematch001_in_ready                        : std_logic;
  signal Kernel_inst_rematch001_in_dvalid                       : std_logic;
  signal Kernel_inst_rematch001_in_last                         : std_logic;
  signal Kernel_inst_rematch001_in_length                       : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch001_in_count                        : std_logic_vector(0 downto 0);
  signal Kernel_inst_rematch001_in_chars_valid                  : std_logic;
  signal Kernel_inst_rematch001_in_chars_ready                  : std_logic;
  signal Kernel_inst_rematch001_in_chars_dvalid                 : std_logic;
  signal Kernel_inst_rematch001_in_chars_last                   : std_logic;
  signal Kernel_inst_rematch001_in_chars                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch001_in_chars_count                  : std_logic_vector(2 downto 0);

  signal Kernel_inst_rematch001_in_unl_valid                    : std_logic;
  signal Kernel_inst_rematch001_in_unl_ready                    : std_logic;
  signal Kernel_inst_rematch001_in_unl_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch001_in_cmd_valid                    : std_logic;
  signal Kernel_inst_rematch001_in_cmd_ready                    : std_logic;
  signal Kernel_inst_rematch001_in_cmd_firstIdx                 : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch001_in_cmd_lastIdx                  : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch001_in_cmd_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch002_in_valid                        : std_logic;
  signal Kernel_inst_rematch002_in_ready                        : std_logic;
  signal Kernel_inst_rematch002_in_dvalid                       : std_logic;
  signal Kernel_inst_rematch002_in_last                         : std_logic;
  signal Kernel_inst_rematch002_in_length                       : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch002_in_count                        : std_logic_vector(0 downto 0);
  signal Kernel_inst_rematch002_in_chars_valid                  : std_logic;
  signal Kernel_inst_rematch002_in_chars_ready                  : std_logic;
  signal Kernel_inst_rematch002_in_chars_dvalid                 : std_logic;
  signal Kernel_inst_rematch002_in_chars_last                   : std_logic;
  signal Kernel_inst_rematch002_in_chars                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch002_in_chars_count                  : std_logic_vector(2 downto 0);

  signal Kernel_inst_rematch002_in_unl_valid                    : std_logic;
  signal Kernel_inst_rematch002_in_unl_ready                    : std_logic;
  signal Kernel_inst_rematch002_in_unl_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch002_in_cmd_valid                    : std_logic;
  signal Kernel_inst_rematch002_in_cmd_ready                    : std_logic;
  signal Kernel_inst_rematch002_in_cmd_firstIdx                 : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch002_in_cmd_lastIdx                  : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch002_in_cmd_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch003_in_valid                        : std_logic;
  signal Kernel_inst_rematch003_in_ready                        : std_logic;
  signal Kernel_inst_rematch003_in_dvalid                       : std_logic;
  signal Kernel_inst_rematch003_in_last                         : std_logic;
  signal Kernel_inst_rematch003_in_length                       : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch003_in_count                        : std_logic_vector(0 downto 0);
  signal Kernel_inst_rematch003_in_chars_valid                  : std_logic;
  signal Kernel_inst_rematch003_in_chars_ready                  : std_logic;
  signal Kernel_inst_rematch003_in_chars_dvalid                 : std_logic;
  signal Kernel_inst_rematch003_in_chars_last                   : std_logic;
  signal Kernel_inst_rematch003_in_chars                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch003_in_chars_count                  : std_logic_vector(2 downto 0);

  signal Kernel_inst_rematch003_in_unl_valid                    : std_logic;
  signal Kernel_inst_rematch003_in_unl_ready                    : std_logic;
  signal Kernel_inst_rematch003_in_unl_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch003_in_cmd_valid                    : std_logic;
  signal Kernel_inst_rematch003_in_cmd_ready                    : std_logic;
  signal Kernel_inst_rematch003_in_cmd_firstIdx                 : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch003_in_cmd_lastIdx                  : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch003_in_cmd_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch004_in_valid                        : std_logic;
  signal Kernel_inst_rematch004_in_ready                        : std_logic;
  signal Kernel_inst_rematch004_in_dvalid                       : std_logic;
  signal Kernel_inst_rematch004_in_last                         : std_logic;
  signal Kernel_inst_rematch004_in_length                       : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch004_in_count                        : std_logic_vector(0 downto 0);
  signal Kernel_inst_rematch004_in_chars_valid                  : std_logic;
  signal Kernel_inst_rematch004_in_chars_ready                  : std_logic;
  signal Kernel_inst_rematch004_in_chars_dvalid                 : std_logic;
  signal Kernel_inst_rematch004_in_chars_last                   : std_logic;
  signal Kernel_inst_rematch004_in_chars                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch004_in_chars_count                  : std_logic_vector(2 downto 0);

  signal Kernel_inst_rematch004_in_unl_valid                    : std_logic;
  signal Kernel_inst_rematch004_in_unl_ready                    : std_logic;
  signal Kernel_inst_rematch004_in_unl_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch004_in_cmd_valid                    : std_logic;
  signal Kernel_inst_rematch004_in_cmd_ready                    : std_logic;
  signal Kernel_inst_rematch004_in_cmd_firstIdx                 : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch004_in_cmd_lastIdx                  : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch004_in_cmd_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch005_in_valid                        : std_logic;
  signal Kernel_inst_rematch005_in_ready                        : std_logic;
  signal Kernel_inst_rematch005_in_dvalid                       : std_logic;
  signal Kernel_inst_rematch005_in_last                         : std_logic;
  signal Kernel_inst_rematch005_in_length                       : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch005_in_count                        : std_logic_vector(0 downto 0);
  signal Kernel_inst_rematch005_in_chars_valid                  : std_logic;
  signal Kernel_inst_rematch005_in_chars_ready                  : std_logic;
  signal Kernel_inst_rematch005_in_chars_dvalid                 : std_logic;
  signal Kernel_inst_rematch005_in_chars_last                   : std_logic;
  signal Kernel_inst_rematch005_in_chars                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch005_in_chars_count                  : std_logic_vector(2 downto 0);

  signal Kernel_inst_rematch005_in_unl_valid                    : std_logic;
  signal Kernel_inst_rematch005_in_unl_ready                    : std_logic;
  signal Kernel_inst_rematch005_in_unl_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch005_in_cmd_valid                    : std_logic;
  signal Kernel_inst_rematch005_in_cmd_ready                    : std_logic;
  signal Kernel_inst_rematch005_in_cmd_firstIdx                 : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch005_in_cmd_lastIdx                  : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch005_in_cmd_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch006_in_valid                        : std_logic;
  signal Kernel_inst_rematch006_in_ready                        : std_logic;
  signal Kernel_inst_rematch006_in_dvalid                       : std_logic;
  signal Kernel_inst_rematch006_in_last                         : std_logic;
  signal Kernel_inst_rematch006_in_length                       : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch006_in_count                        : std_logic_vector(0 downto 0);
  signal Kernel_inst_rematch006_in_chars_valid                  : std_logic;
  signal Kernel_inst_rematch006_in_chars_ready                  : std_logic;
  signal Kernel_inst_rematch006_in_chars_dvalid                 : std_logic;
  signal Kernel_inst_rematch006_in_chars_last                   : std_logic;
  signal Kernel_inst_rematch006_in_chars                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch006_in_chars_count                  : std_logic_vector(2 downto 0);

  signal Kernel_inst_rematch006_in_unl_valid                    : std_logic;
  signal Kernel_inst_rematch006_in_unl_ready                    : std_logic;
  signal Kernel_inst_rematch006_in_unl_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch006_in_cmd_valid                    : std_logic;
  signal Kernel_inst_rematch006_in_cmd_ready                    : std_logic;
  signal Kernel_inst_rematch006_in_cmd_firstIdx                 : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch006_in_cmd_lastIdx                  : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch006_in_cmd_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch007_in_valid                        : std_logic;
  signal Kernel_inst_rematch007_in_ready                        : std_logic;
  signal Kernel_inst_rematch007_in_dvalid                       : std_logic;
  signal Kernel_inst_rematch007_in_last                         : std_logic;
  signal Kernel_inst_rematch007_in_length                       : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch007_in_count                        : std_logic_vector(0 downto 0);
  signal Kernel_inst_rematch007_in_chars_valid                  : std_logic;
  signal Kernel_inst_rematch007_in_chars_ready                  : std_logic;
  signal Kernel_inst_rematch007_in_chars_dvalid                 : std_logic;
  signal Kernel_inst_rematch007_in_chars_last                   : std_logic;
  signal Kernel_inst_rematch007_in_chars                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch007_in_chars_count                  : std_logic_vector(2 downto 0);

  signal Kernel_inst_rematch007_in_unl_valid                    : std_logic;
  signal Kernel_inst_rematch007_in_unl_ready                    : std_logic;
  signal Kernel_inst_rematch007_in_unl_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch007_in_cmd_valid                    : std_logic;
  signal Kernel_inst_rematch007_in_cmd_ready                    : std_logic;
  signal Kernel_inst_rematch007_in_cmd_firstIdx                 : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch007_in_cmd_lastIdx                  : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch007_in_cmd_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch008_in_valid                        : std_logic;
  signal Kernel_inst_rematch008_in_ready                        : std_logic;
  signal Kernel_inst_rematch008_in_dvalid                       : std_logic;
  signal Kernel_inst_rematch008_in_last                         : std_logic;
  signal Kernel_inst_rematch008_in_length                       : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch008_in_count                        : std_logic_vector(0 downto 0);
  signal Kernel_inst_rematch008_in_chars_valid                  : std_logic;
  signal Kernel_inst_rematch008_in_chars_ready                  : std_logic;
  signal Kernel_inst_rematch008_in_chars_dvalid                 : std_logic;
  signal Kernel_inst_rematch008_in_chars_last                   : std_logic;
  signal Kernel_inst_rematch008_in_chars                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch008_in_chars_count                  : std_logic_vector(2 downto 0);

  signal Kernel_inst_rematch008_in_unl_valid                    : std_logic;
  signal Kernel_inst_rematch008_in_unl_ready                    : std_logic;
  signal Kernel_inst_rematch008_in_unl_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch008_in_cmd_valid                    : std_logic;
  signal Kernel_inst_rematch008_in_cmd_ready                    : std_logic;
  signal Kernel_inst_rematch008_in_cmd_firstIdx                 : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch008_in_cmd_lastIdx                  : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch008_in_cmd_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch009_in_valid                        : std_logic;
  signal Kernel_inst_rematch009_in_ready                        : std_logic;
  signal Kernel_inst_rematch009_in_dvalid                       : std_logic;
  signal Kernel_inst_rematch009_in_last                         : std_logic;
  signal Kernel_inst_rematch009_in_length                       : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch009_in_count                        : std_logic_vector(0 downto 0);
  signal Kernel_inst_rematch009_in_chars_valid                  : std_logic;
  signal Kernel_inst_rematch009_in_chars_ready                  : std_logic;
  signal Kernel_inst_rematch009_in_chars_dvalid                 : std_logic;
  signal Kernel_inst_rematch009_in_chars_last                   : std_logic;
  signal Kernel_inst_rematch009_in_chars                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch009_in_chars_count                  : std_logic_vector(2 downto 0);

  signal Kernel_inst_rematch009_in_unl_valid                    : std_logic;
  signal Kernel_inst_rematch009_in_unl_ready                    : std_logic;
  signal Kernel_inst_rematch009_in_unl_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch009_in_cmd_valid                    : std_logic;
  signal Kernel_inst_rematch009_in_cmd_ready                    : std_logic;
  signal Kernel_inst_rematch009_in_cmd_firstIdx                 : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch009_in_cmd_lastIdx                  : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch009_in_cmd_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch010_in_valid                        : std_logic;
  signal Kernel_inst_rematch010_in_ready                        : std_logic;
  signal Kernel_inst_rematch010_in_dvalid                       : std_logic;
  signal Kernel_inst_rematch010_in_last                         : std_logic;
  signal Kernel_inst_rematch010_in_length                       : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch010_in_count                        : std_logic_vector(0 downto 0);
  signal Kernel_inst_rematch010_in_chars_valid                  : std_logic;
  signal Kernel_inst_rematch010_in_chars_ready                  : std_logic;
  signal Kernel_inst_rematch010_in_chars_dvalid                 : std_logic;
  signal Kernel_inst_rematch010_in_chars_last                   : std_logic;
  signal Kernel_inst_rematch010_in_chars                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch010_in_chars_count                  : std_logic_vector(2 downto 0);

  signal Kernel_inst_rematch010_in_unl_valid                    : std_logic;
  signal Kernel_inst_rematch010_in_unl_ready                    : std_logic;
  signal Kernel_inst_rematch010_in_unl_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch010_in_cmd_valid                    : std_logic;
  signal Kernel_inst_rematch010_in_cmd_ready                    : std_logic;
  signal Kernel_inst_rematch010_in_cmd_firstIdx                 : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch010_in_cmd_lastIdx                  : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch010_in_cmd_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch011_in_valid                        : std_logic;
  signal Kernel_inst_rematch011_in_ready                        : std_logic;
  signal Kernel_inst_rematch011_in_dvalid                       : std_logic;
  signal Kernel_inst_rematch011_in_last                         : std_logic;
  signal Kernel_inst_rematch011_in_length                       : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch011_in_count                        : std_logic_vector(0 downto 0);
  signal Kernel_inst_rematch011_in_chars_valid                  : std_logic;
  signal Kernel_inst_rematch011_in_chars_ready                  : std_logic;
  signal Kernel_inst_rematch011_in_chars_dvalid                 : std_logic;
  signal Kernel_inst_rematch011_in_chars_last                   : std_logic;
  signal Kernel_inst_rematch011_in_chars                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch011_in_chars_count                  : std_logic_vector(2 downto 0);

  signal Kernel_inst_rematch011_in_unl_valid                    : std_logic;
  signal Kernel_inst_rematch011_in_unl_ready                    : std_logic;
  signal Kernel_inst_rematch011_in_unl_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch011_in_cmd_valid                    : std_logic;
  signal Kernel_inst_rematch011_in_cmd_ready                    : std_logic;
  signal Kernel_inst_rematch011_in_cmd_firstIdx                 : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch011_in_cmd_lastIdx                  : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch011_in_cmd_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch012_in_valid                        : std_logic;
  signal Kernel_inst_rematch012_in_ready                        : std_logic;
  signal Kernel_inst_rematch012_in_dvalid                       : std_logic;
  signal Kernel_inst_rematch012_in_last                         : std_logic;
  signal Kernel_inst_rematch012_in_length                       : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch012_in_count                        : std_logic_vector(0 downto 0);
  signal Kernel_inst_rematch012_in_chars_valid                  : std_logic;
  signal Kernel_inst_rematch012_in_chars_ready                  : std_logic;
  signal Kernel_inst_rematch012_in_chars_dvalid                 : std_logic;
  signal Kernel_inst_rematch012_in_chars_last                   : std_logic;
  signal Kernel_inst_rematch012_in_chars                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch012_in_chars_count                  : std_logic_vector(2 downto 0);

  signal Kernel_inst_rematch012_in_unl_valid                    : std_logic;
  signal Kernel_inst_rematch012_in_unl_ready                    : std_logic;
  signal Kernel_inst_rematch012_in_unl_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch012_in_cmd_valid                    : std_logic;
  signal Kernel_inst_rematch012_in_cmd_ready                    : std_logic;
  signal Kernel_inst_rematch012_in_cmd_firstIdx                 : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch012_in_cmd_lastIdx                  : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch012_in_cmd_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch013_in_valid                        : std_logic;
  signal Kernel_inst_rematch013_in_ready                        : std_logic;
  signal Kernel_inst_rematch013_in_dvalid                       : std_logic;
  signal Kernel_inst_rematch013_in_last                         : std_logic;
  signal Kernel_inst_rematch013_in_length                       : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch013_in_count                        : std_logic_vector(0 downto 0);
  signal Kernel_inst_rematch013_in_chars_valid                  : std_logic;
  signal Kernel_inst_rematch013_in_chars_ready                  : std_logic;
  signal Kernel_inst_rematch013_in_chars_dvalid                 : std_logic;
  signal Kernel_inst_rematch013_in_chars_last                   : std_logic;
  signal Kernel_inst_rematch013_in_chars                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch013_in_chars_count                  : std_logic_vector(2 downto 0);

  signal Kernel_inst_rematch013_in_unl_valid                    : std_logic;
  signal Kernel_inst_rematch013_in_unl_ready                    : std_logic;
  signal Kernel_inst_rematch013_in_unl_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch013_in_cmd_valid                    : std_logic;
  signal Kernel_inst_rematch013_in_cmd_ready                    : std_logic;
  signal Kernel_inst_rematch013_in_cmd_firstIdx                 : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch013_in_cmd_lastIdx                  : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch013_in_cmd_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch014_in_valid                        : std_logic;
  signal Kernel_inst_rematch014_in_ready                        : std_logic;
  signal Kernel_inst_rematch014_in_dvalid                       : std_logic;
  signal Kernel_inst_rematch014_in_last                         : std_logic;
  signal Kernel_inst_rematch014_in_length                       : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch014_in_count                        : std_logic_vector(0 downto 0);
  signal Kernel_inst_rematch014_in_chars_valid                  : std_logic;
  signal Kernel_inst_rematch014_in_chars_ready                  : std_logic;
  signal Kernel_inst_rematch014_in_chars_dvalid                 : std_logic;
  signal Kernel_inst_rematch014_in_chars_last                   : std_logic;
  signal Kernel_inst_rematch014_in_chars                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch014_in_chars_count                  : std_logic_vector(2 downto 0);

  signal Kernel_inst_rematch014_in_unl_valid                    : std_logic;
  signal Kernel_inst_rematch014_in_unl_ready                    : std_logic;
  signal Kernel_inst_rematch014_in_unl_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch014_in_cmd_valid                    : std_logic;
  signal Kernel_inst_rematch014_in_cmd_ready                    : std_logic;
  signal Kernel_inst_rematch014_in_cmd_firstIdx                 : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch014_in_cmd_lastIdx                  : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch014_in_cmd_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch015_in_valid                        : std_logic;
  signal Kernel_inst_rematch015_in_ready                        : std_logic;
  signal Kernel_inst_rematch015_in_dvalid                       : std_logic;
  signal Kernel_inst_rematch015_in_last                         : std_logic;
  signal Kernel_inst_rematch015_in_length                       : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch015_in_count                        : std_logic_vector(0 downto 0);
  signal Kernel_inst_rematch015_in_chars_valid                  : std_logic;
  signal Kernel_inst_rematch015_in_chars_ready                  : std_logic;
  signal Kernel_inst_rematch015_in_chars_dvalid                 : std_logic;
  signal Kernel_inst_rematch015_in_chars_last                   : std_logic;
  signal Kernel_inst_rematch015_in_chars                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch015_in_chars_count                  : std_logic_vector(2 downto 0);

  signal Kernel_inst_rematch015_in_unl_valid                    : std_logic;
  signal Kernel_inst_rematch015_in_unl_ready                    : std_logic;
  signal Kernel_inst_rematch015_in_unl_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch015_in_cmd_valid                    : std_logic;
  signal Kernel_inst_rematch015_in_cmd_ready                    : std_logic;
  signal Kernel_inst_rematch015_in_cmd_firstIdx                 : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch015_in_cmd_lastIdx                  : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch015_in_cmd_tag                      : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch000_taxi_out_valid                  : std_logic;
  signal Kernel_inst_rematch000_taxi_out_ready                  : std_logic;
  signal Kernel_inst_rematch000_taxi_out_dvalid                 : std_logic;
  signal Kernel_inst_rematch000_taxi_out_last                   : std_logic;
  signal Kernel_inst_rematch000_taxi_out                        : std_logic_vector(31 downto 0);

  signal Kernel_inst_rematch000_taxi_out_unl_valid              : std_logic;
  signal Kernel_inst_rematch000_taxi_out_unl_ready              : std_logic;
  signal Kernel_inst_rematch000_taxi_out_unl_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch000_taxi_out_cmd_valid              : std_logic;
  signal Kernel_inst_rematch000_taxi_out_cmd_ready              : std_logic;
  signal Kernel_inst_rematch000_taxi_out_cmd_firstIdx           : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch000_taxi_out_cmd_lastIdx            : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch000_taxi_out_cmd_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch001_taxi_out_valid                  : std_logic;
  signal Kernel_inst_rematch001_taxi_out_ready                  : std_logic;
  signal Kernel_inst_rematch001_taxi_out_dvalid                 : std_logic;
  signal Kernel_inst_rematch001_taxi_out_last                   : std_logic;
  signal Kernel_inst_rematch001_taxi_out                        : std_logic_vector(31 downto 0);

  signal Kernel_inst_rematch001_taxi_out_unl_valid              : std_logic;
  signal Kernel_inst_rematch001_taxi_out_unl_ready              : std_logic;
  signal Kernel_inst_rematch001_taxi_out_unl_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch001_taxi_out_cmd_valid              : std_logic;
  signal Kernel_inst_rematch001_taxi_out_cmd_ready              : std_logic;
  signal Kernel_inst_rematch001_taxi_out_cmd_firstIdx           : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch001_taxi_out_cmd_lastIdx            : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch001_taxi_out_cmd_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch002_taxi_out_valid                  : std_logic;
  signal Kernel_inst_rematch002_taxi_out_ready                  : std_logic;
  signal Kernel_inst_rematch002_taxi_out_dvalid                 : std_logic;
  signal Kernel_inst_rematch002_taxi_out_last                   : std_logic;
  signal Kernel_inst_rematch002_taxi_out                        : std_logic_vector(31 downto 0);

  signal Kernel_inst_rematch002_taxi_out_unl_valid              : std_logic;
  signal Kernel_inst_rematch002_taxi_out_unl_ready              : std_logic;
  signal Kernel_inst_rematch002_taxi_out_unl_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch002_taxi_out_cmd_valid              : std_logic;
  signal Kernel_inst_rematch002_taxi_out_cmd_ready              : std_logic;
  signal Kernel_inst_rematch002_taxi_out_cmd_firstIdx           : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch002_taxi_out_cmd_lastIdx            : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch002_taxi_out_cmd_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch003_taxi_out_valid                  : std_logic;
  signal Kernel_inst_rematch003_taxi_out_ready                  : std_logic;
  signal Kernel_inst_rematch003_taxi_out_dvalid                 : std_logic;
  signal Kernel_inst_rematch003_taxi_out_last                   : std_logic;
  signal Kernel_inst_rematch003_taxi_out                        : std_logic_vector(31 downto 0);

  signal Kernel_inst_rematch003_taxi_out_unl_valid              : std_logic;
  signal Kernel_inst_rematch003_taxi_out_unl_ready              : std_logic;
  signal Kernel_inst_rematch003_taxi_out_unl_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch003_taxi_out_cmd_valid              : std_logic;
  signal Kernel_inst_rematch003_taxi_out_cmd_ready              : std_logic;
  signal Kernel_inst_rematch003_taxi_out_cmd_firstIdx           : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch003_taxi_out_cmd_lastIdx            : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch003_taxi_out_cmd_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch004_taxi_out_valid                  : std_logic;
  signal Kernel_inst_rematch004_taxi_out_ready                  : std_logic;
  signal Kernel_inst_rematch004_taxi_out_dvalid                 : std_logic;
  signal Kernel_inst_rematch004_taxi_out_last                   : std_logic;
  signal Kernel_inst_rematch004_taxi_out                        : std_logic_vector(31 downto 0);

  signal Kernel_inst_rematch004_taxi_out_unl_valid              : std_logic;
  signal Kernel_inst_rematch004_taxi_out_unl_ready              : std_logic;
  signal Kernel_inst_rematch004_taxi_out_unl_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch004_taxi_out_cmd_valid              : std_logic;
  signal Kernel_inst_rematch004_taxi_out_cmd_ready              : std_logic;
  signal Kernel_inst_rematch004_taxi_out_cmd_firstIdx           : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch004_taxi_out_cmd_lastIdx            : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch004_taxi_out_cmd_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch005_taxi_out_valid                  : std_logic;
  signal Kernel_inst_rematch005_taxi_out_ready                  : std_logic;
  signal Kernel_inst_rematch005_taxi_out_dvalid                 : std_logic;
  signal Kernel_inst_rematch005_taxi_out_last                   : std_logic;
  signal Kernel_inst_rematch005_taxi_out                        : std_logic_vector(31 downto 0);

  signal Kernel_inst_rematch005_taxi_out_unl_valid              : std_logic;
  signal Kernel_inst_rematch005_taxi_out_unl_ready              : std_logic;
  signal Kernel_inst_rematch005_taxi_out_unl_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch005_taxi_out_cmd_valid              : std_logic;
  signal Kernel_inst_rematch005_taxi_out_cmd_ready              : std_logic;
  signal Kernel_inst_rematch005_taxi_out_cmd_firstIdx           : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch005_taxi_out_cmd_lastIdx            : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch005_taxi_out_cmd_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch006_taxi_out_valid                  : std_logic;
  signal Kernel_inst_rematch006_taxi_out_ready                  : std_logic;
  signal Kernel_inst_rematch006_taxi_out_dvalid                 : std_logic;
  signal Kernel_inst_rematch006_taxi_out_last                   : std_logic;
  signal Kernel_inst_rematch006_taxi_out                        : std_logic_vector(31 downto 0);

  signal Kernel_inst_rematch006_taxi_out_unl_valid              : std_logic;
  signal Kernel_inst_rematch006_taxi_out_unl_ready              : std_logic;
  signal Kernel_inst_rematch006_taxi_out_unl_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch006_taxi_out_cmd_valid              : std_logic;
  signal Kernel_inst_rematch006_taxi_out_cmd_ready              : std_logic;
  signal Kernel_inst_rematch006_taxi_out_cmd_firstIdx           : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch006_taxi_out_cmd_lastIdx            : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch006_taxi_out_cmd_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch007_taxi_out_valid                  : std_logic;
  signal Kernel_inst_rematch007_taxi_out_ready                  : std_logic;
  signal Kernel_inst_rematch007_taxi_out_dvalid                 : std_logic;
  signal Kernel_inst_rematch007_taxi_out_last                   : std_logic;
  signal Kernel_inst_rematch007_taxi_out                        : std_logic_vector(31 downto 0);

  signal Kernel_inst_rematch007_taxi_out_unl_valid              : std_logic;
  signal Kernel_inst_rematch007_taxi_out_unl_ready              : std_logic;
  signal Kernel_inst_rematch007_taxi_out_unl_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch007_taxi_out_cmd_valid              : std_logic;
  signal Kernel_inst_rematch007_taxi_out_cmd_ready              : std_logic;
  signal Kernel_inst_rematch007_taxi_out_cmd_firstIdx           : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch007_taxi_out_cmd_lastIdx            : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch007_taxi_out_cmd_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch008_taxi_out_valid                  : std_logic;
  signal Kernel_inst_rematch008_taxi_out_ready                  : std_logic;
  signal Kernel_inst_rematch008_taxi_out_dvalid                 : std_logic;
  signal Kernel_inst_rematch008_taxi_out_last                   : std_logic;
  signal Kernel_inst_rematch008_taxi_out                        : std_logic_vector(31 downto 0);

  signal Kernel_inst_rematch008_taxi_out_unl_valid              : std_logic;
  signal Kernel_inst_rematch008_taxi_out_unl_ready              : std_logic;
  signal Kernel_inst_rematch008_taxi_out_unl_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch008_taxi_out_cmd_valid              : std_logic;
  signal Kernel_inst_rematch008_taxi_out_cmd_ready              : std_logic;
  signal Kernel_inst_rematch008_taxi_out_cmd_firstIdx           : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch008_taxi_out_cmd_lastIdx            : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch008_taxi_out_cmd_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch009_taxi_out_valid                  : std_logic;
  signal Kernel_inst_rematch009_taxi_out_ready                  : std_logic;
  signal Kernel_inst_rematch009_taxi_out_dvalid                 : std_logic;
  signal Kernel_inst_rematch009_taxi_out_last                   : std_logic;
  signal Kernel_inst_rematch009_taxi_out                        : std_logic_vector(31 downto 0);

  signal Kernel_inst_rematch009_taxi_out_unl_valid              : std_logic;
  signal Kernel_inst_rematch009_taxi_out_unl_ready              : std_logic;
  signal Kernel_inst_rematch009_taxi_out_unl_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch009_taxi_out_cmd_valid              : std_logic;
  signal Kernel_inst_rematch009_taxi_out_cmd_ready              : std_logic;
  signal Kernel_inst_rematch009_taxi_out_cmd_firstIdx           : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch009_taxi_out_cmd_lastIdx            : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch009_taxi_out_cmd_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch010_taxi_out_valid                  : std_logic;
  signal Kernel_inst_rematch010_taxi_out_ready                  : std_logic;
  signal Kernel_inst_rematch010_taxi_out_dvalid                 : std_logic;
  signal Kernel_inst_rematch010_taxi_out_last                   : std_logic;
  signal Kernel_inst_rematch010_taxi_out                        : std_logic_vector(31 downto 0);

  signal Kernel_inst_rematch010_taxi_out_unl_valid              : std_logic;
  signal Kernel_inst_rematch010_taxi_out_unl_ready              : std_logic;
  signal Kernel_inst_rematch010_taxi_out_unl_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch010_taxi_out_cmd_valid              : std_logic;
  signal Kernel_inst_rematch010_taxi_out_cmd_ready              : std_logic;
  signal Kernel_inst_rematch010_taxi_out_cmd_firstIdx           : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch010_taxi_out_cmd_lastIdx            : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch010_taxi_out_cmd_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch011_taxi_out_valid                  : std_logic;
  signal Kernel_inst_rematch011_taxi_out_ready                  : std_logic;
  signal Kernel_inst_rematch011_taxi_out_dvalid                 : std_logic;
  signal Kernel_inst_rematch011_taxi_out_last                   : std_logic;
  signal Kernel_inst_rematch011_taxi_out                        : std_logic_vector(31 downto 0);

  signal Kernel_inst_rematch011_taxi_out_unl_valid              : std_logic;
  signal Kernel_inst_rematch011_taxi_out_unl_ready              : std_logic;
  signal Kernel_inst_rematch011_taxi_out_unl_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch011_taxi_out_cmd_valid              : std_logic;
  signal Kernel_inst_rematch011_taxi_out_cmd_ready              : std_logic;
  signal Kernel_inst_rematch011_taxi_out_cmd_firstIdx           : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch011_taxi_out_cmd_lastIdx            : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch011_taxi_out_cmd_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch012_taxi_out_valid                  : std_logic;
  signal Kernel_inst_rematch012_taxi_out_ready                  : std_logic;
  signal Kernel_inst_rematch012_taxi_out_dvalid                 : std_logic;
  signal Kernel_inst_rematch012_taxi_out_last                   : std_logic;
  signal Kernel_inst_rematch012_taxi_out                        : std_logic_vector(31 downto 0);

  signal Kernel_inst_rematch012_taxi_out_unl_valid              : std_logic;
  signal Kernel_inst_rematch012_taxi_out_unl_ready              : std_logic;
  signal Kernel_inst_rematch012_taxi_out_unl_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch012_taxi_out_cmd_valid              : std_logic;
  signal Kernel_inst_rematch012_taxi_out_cmd_ready              : std_logic;
  signal Kernel_inst_rematch012_taxi_out_cmd_firstIdx           : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch012_taxi_out_cmd_lastIdx            : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch012_taxi_out_cmd_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch013_taxi_out_valid                  : std_logic;
  signal Kernel_inst_rematch013_taxi_out_ready                  : std_logic;
  signal Kernel_inst_rematch013_taxi_out_dvalid                 : std_logic;
  signal Kernel_inst_rematch013_taxi_out_last                   : std_logic;
  signal Kernel_inst_rematch013_taxi_out                        : std_logic_vector(31 downto 0);

  signal Kernel_inst_rematch013_taxi_out_unl_valid              : std_logic;
  signal Kernel_inst_rematch013_taxi_out_unl_ready              : std_logic;
  signal Kernel_inst_rematch013_taxi_out_unl_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch013_taxi_out_cmd_valid              : std_logic;
  signal Kernel_inst_rematch013_taxi_out_cmd_ready              : std_logic;
  signal Kernel_inst_rematch013_taxi_out_cmd_firstIdx           : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch013_taxi_out_cmd_lastIdx            : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch013_taxi_out_cmd_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch014_taxi_out_valid                  : std_logic;
  signal Kernel_inst_rematch014_taxi_out_ready                  : std_logic;
  signal Kernel_inst_rematch014_taxi_out_dvalid                 : std_logic;
  signal Kernel_inst_rematch014_taxi_out_last                   : std_logic;
  signal Kernel_inst_rematch014_taxi_out                        : std_logic_vector(31 downto 0);

  signal Kernel_inst_rematch014_taxi_out_unl_valid              : std_logic;
  signal Kernel_inst_rematch014_taxi_out_unl_ready              : std_logic;
  signal Kernel_inst_rematch014_taxi_out_unl_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch014_taxi_out_cmd_valid              : std_logic;
  signal Kernel_inst_rematch014_taxi_out_cmd_ready              : std_logic;
  signal Kernel_inst_rematch014_taxi_out_cmd_firstIdx           : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch014_taxi_out_cmd_lastIdx            : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch014_taxi_out_cmd_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch015_taxi_out_valid                  : std_logic;
  signal Kernel_inst_rematch015_taxi_out_ready                  : std_logic;
  signal Kernel_inst_rematch015_taxi_out_dvalid                 : std_logic;
  signal Kernel_inst_rematch015_taxi_out_last                   : std_logic;
  signal Kernel_inst_rematch015_taxi_out                        : std_logic_vector(31 downto 0);

  signal Kernel_inst_rematch015_taxi_out_unl_valid              : std_logic;
  signal Kernel_inst_rematch015_taxi_out_unl_ready              : std_logic;
  signal Kernel_inst_rematch015_taxi_out_unl_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_rematch015_taxi_out_cmd_valid              : std_logic;
  signal Kernel_inst_rematch015_taxi_out_cmd_ready              : std_logic;
  signal Kernel_inst_rematch015_taxi_out_cmd_firstIdx           : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch015_taxi_out_cmd_lastIdx            : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch015_taxi_out_cmd_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_start                                      : std_logic;
  signal Kernel_inst_stop                                       : std_logic;
  signal Kernel_inst_reset                                      : std_logic;
  signal Kernel_inst_idle                                       : std_logic;
  signal Kernel_inst_busy                                       : std_logic;
  signal Kernel_inst_done                                       : std_logic;
  signal Kernel_inst_result                                     : std_logic_vector(63 downto 0);
  signal Kernel_inst_rematch000_firstidx                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch000_lastidx                         : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch001_firstidx                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch001_lastidx                         : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch002_firstidx                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch002_lastidx                         : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch003_firstidx                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch003_lastidx                         : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch004_firstidx                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch004_lastidx                         : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch005_firstidx                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch005_lastidx                         : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch006_firstidx                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch006_lastidx                         : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch007_firstidx                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch007_lastidx                         : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch008_firstidx                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch008_lastidx                         : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch009_firstidx                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch009_lastidx                         : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch010_firstidx                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch010_lastidx                         : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch011_firstidx                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch011_lastidx                         : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch012_firstidx                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch012_lastidx                         : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch013_firstidx                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch013_lastidx                         : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch014_firstidx                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch014_lastidx                         : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch015_firstidx                        : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch015_lastidx                         : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch000_taxi_firstidx                   : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch000_taxi_lastidx                    : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch001_taxi_firstidx                   : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch001_taxi_lastidx                    : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch002_taxi_firstidx                   : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch002_taxi_lastidx                    : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch003_taxi_firstidx                   : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch003_taxi_lastidx                    : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch004_taxi_firstidx                   : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch004_taxi_lastidx                    : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch005_taxi_firstidx                   : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch005_taxi_lastidx                    : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch006_taxi_firstidx                   : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch006_taxi_lastidx                    : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch007_taxi_firstidx                   : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch007_taxi_lastidx                    : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch008_taxi_firstidx                   : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch008_taxi_lastidx                    : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch009_taxi_firstidx                   : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch009_taxi_lastidx                    : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch010_taxi_firstidx                   : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch010_taxi_lastidx                    : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch011_taxi_firstidx                   : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch011_taxi_lastidx                    : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch012_taxi_firstidx                   : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch012_taxi_lastidx                    : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch013_taxi_firstidx                   : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch013_taxi_lastidx                    : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch014_taxi_firstidx                   : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch014_taxi_lastidx                    : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch015_taxi_firstidx                   : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch015_taxi_lastidx                    : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch000_taxi_count                      : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch000_errors                          : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch001_taxi_count                      : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch001_errors                          : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch002_taxi_count                      : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch002_errors                          : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch003_taxi_count                      : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch003_errors                          : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch004_taxi_count                      : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch004_errors                          : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch005_taxi_count                      : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch005_errors                          : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch006_taxi_count                      : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch006_errors                          : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch007_taxi_count                      : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch007_errors                          : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch008_taxi_count                      : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch008_errors                          : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch009_taxi_count                      : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch009_errors                          : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch010_taxi_count                      : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch010_errors                          : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch011_taxi_count                      : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch011_errors                          : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch012_taxi_count                      : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch012_errors                          : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch013_taxi_count                      : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch013_errors                          : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch014_taxi_count                      : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch014_errors                          : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch015_taxi_count                      : std_logic_vector(31 downto 0);
  signal Kernel_inst_rematch015_errors                          : std_logic_vector(31 downto 0);
  signal mmio_inst_f_start_data                                 : std_logic;
  signal mmio_inst_f_stop_data                                  : std_logic;
  signal mmio_inst_f_reset_data                                 : std_logic;
  signal mmio_inst_f_idle_write_data                            : std_logic;
  signal mmio_inst_f_busy_write_data                            : std_logic;
  signal mmio_inst_f_done_write_data                            : std_logic;
  signal mmio_inst_f_result_write_data                          : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch000_firstidx_data                   : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch000_lastidx_data                    : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch001_firstidx_data                   : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch001_lastidx_data                    : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch002_firstidx_data                   : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch002_lastidx_data                    : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch003_firstidx_data                   : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch003_lastidx_data                    : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch004_firstidx_data                   : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch004_lastidx_data                    : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch005_firstidx_data                   : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch005_lastidx_data                    : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch006_firstidx_data                   : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch006_lastidx_data                    : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch007_firstidx_data                   : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch007_lastidx_data                    : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch008_firstidx_data                   : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch008_lastidx_data                    : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch009_firstidx_data                   : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch009_lastidx_data                    : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch010_firstidx_data                   : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch010_lastidx_data                    : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch011_firstidx_data                   : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch011_lastidx_data                    : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch012_firstidx_data                   : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch012_lastidx_data                    : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch013_firstidx_data                   : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch013_lastidx_data                    : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch014_firstidx_data                   : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch014_lastidx_data                    : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch015_firstidx_data                   : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch015_lastidx_data                    : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch000_taxi_firstidx_data              : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch000_taxi_lastidx_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch001_taxi_firstidx_data              : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch001_taxi_lastidx_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch002_taxi_firstidx_data              : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch002_taxi_lastidx_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch003_taxi_firstidx_data              : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch003_taxi_lastidx_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch004_taxi_firstidx_data              : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch004_taxi_lastidx_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch005_taxi_firstidx_data              : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch005_taxi_lastidx_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch006_taxi_firstidx_data              : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch006_taxi_lastidx_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch007_taxi_firstidx_data              : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch007_taxi_lastidx_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch008_taxi_firstidx_data              : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch008_taxi_lastidx_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch009_taxi_firstidx_data              : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch009_taxi_lastidx_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch010_taxi_firstidx_data              : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch010_taxi_lastidx_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch011_taxi_firstidx_data              : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch011_taxi_lastidx_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch012_taxi_firstidx_data              : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch012_taxi_lastidx_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch013_taxi_firstidx_data              : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch013_taxi_lastidx_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch014_taxi_firstidx_data              : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch014_taxi_lastidx_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch015_taxi_firstidx_data              : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch015_taxi_lastidx_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch000_in_offsets_data                 : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch000_in_values_data                  : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch001_in_offsets_data                 : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch001_in_values_data                  : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch002_in_offsets_data                 : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch002_in_values_data                  : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch003_in_offsets_data                 : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch003_in_values_data                  : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch004_in_offsets_data                 : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch004_in_values_data                  : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch005_in_offsets_data                 : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch005_in_values_data                  : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch006_in_offsets_data                 : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch006_in_values_data                  : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch007_in_offsets_data                 : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch007_in_values_data                  : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch008_in_offsets_data                 : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch008_in_values_data                  : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch009_in_offsets_data                 : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch009_in_values_data                  : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch010_in_offsets_data                 : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch010_in_values_data                  : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch011_in_offsets_data                 : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch011_in_values_data                  : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch012_in_offsets_data                 : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch012_in_values_data                  : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch013_in_offsets_data                 : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch013_in_values_data                  : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch014_in_offsets_data                 : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch014_in_values_data                  : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch015_in_offsets_data                 : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch015_in_values_data                  : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch000_taxi_out_values_data            : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch001_taxi_out_values_data            : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch002_taxi_out_values_data            : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch003_taxi_out_values_data            : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch004_taxi_out_values_data            : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch005_taxi_out_values_data            : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch006_taxi_out_values_data            : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch007_taxi_out_values_data            : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch008_taxi_out_values_data            : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch009_taxi_out_values_data            : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch010_taxi_out_values_data            : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch011_taxi_out_values_data            : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch012_taxi_out_values_data            : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch013_taxi_out_values_data            : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch014_taxi_out_values_data            : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch015_taxi_out_values_data            : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rematch000_taxi_count_write_data           : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch000_errors_write_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch001_taxi_count_write_data           : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch001_errors_write_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch002_taxi_count_write_data           : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch002_errors_write_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch003_taxi_count_write_data           : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch003_errors_write_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch004_taxi_count_write_data           : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch004_errors_write_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch005_taxi_count_write_data           : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch005_errors_write_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch006_taxi_count_write_data           : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch006_errors_write_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch007_taxi_count_write_data           : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch007_errors_write_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch008_taxi_count_write_data           : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch008_errors_write_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch009_taxi_count_write_data           : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch009_errors_write_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch010_taxi_count_write_data           : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch010_errors_write_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch011_taxi_count_write_data           : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch011_errors_write_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch012_taxi_count_write_data           : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch012_errors_write_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch013_taxi_count_write_data           : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch013_errors_write_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch014_taxi_count_write_data           : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch014_errors_write_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch015_taxi_count_write_data           : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rematch015_errors_write_data               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_Profile_enable_data                        : std_logic;
  signal mmio_inst_f_Profile_clear_data                         : std_logic;
  signal mmio_inst_mmio_awvalid                                 : std_logic;
  signal mmio_inst_mmio_awready                                 : std_logic;
  signal mmio_inst_mmio_awaddr                                  : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_wvalid                                  : std_logic;
  signal mmio_inst_mmio_wready                                  : std_logic;
  signal mmio_inst_mmio_wdata                                   : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_wstrb                                   : std_logic_vector(3 downto 0);
  signal mmio_inst_mmio_bvalid                                  : std_logic;
  signal mmio_inst_mmio_bready                                  : std_logic;
  signal mmio_inst_mmio_bresp                                   : std_logic_vector(1 downto 0);
  signal mmio_inst_mmio_arvalid                                 : std_logic;
  signal mmio_inst_mmio_arready                                 : std_logic;
  signal mmio_inst_mmio_araddr                                  : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_rvalid                                  : std_logic;
  signal mmio_inst_mmio_rready                                  : std_logic;
  signal mmio_inst_mmio_rdata                                   : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_rresp                                   : std_logic_vector(1 downto 0);

  signal rematch000_in_cmd_accm_inst_kernel_cmd_valid           : std_logic;
  signal rematch000_in_cmd_accm_inst_kernel_cmd_ready           : std_logic;
  signal rematch000_in_cmd_accm_inst_kernel_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch000_in_cmd_accm_inst_kernel_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch000_in_cmd_accm_inst_kernel_cmd_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch000_in_cmd_accm_inst_nucleus_cmd_valid          : std_logic;
  signal rematch000_in_cmd_accm_inst_nucleus_cmd_ready          : std_logic;
  signal rematch000_in_cmd_accm_inst_nucleus_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch000_in_cmd_accm_inst_nucleus_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch000_in_cmd_accm_inst_nucleus_cmd_ctrl           : std_logic_vector(2*REMATCH000_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch000_in_cmd_accm_inst_nucleus_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch001_in_cmd_accm_inst_kernel_cmd_valid           : std_logic;
  signal rematch001_in_cmd_accm_inst_kernel_cmd_ready           : std_logic;
  signal rematch001_in_cmd_accm_inst_kernel_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch001_in_cmd_accm_inst_kernel_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch001_in_cmd_accm_inst_kernel_cmd_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch001_in_cmd_accm_inst_nucleus_cmd_valid          : std_logic;
  signal rematch001_in_cmd_accm_inst_nucleus_cmd_ready          : std_logic;
  signal rematch001_in_cmd_accm_inst_nucleus_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch001_in_cmd_accm_inst_nucleus_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch001_in_cmd_accm_inst_nucleus_cmd_ctrl           : std_logic_vector(2*REMATCH001_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch001_in_cmd_accm_inst_nucleus_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch002_in_cmd_accm_inst_kernel_cmd_valid           : std_logic;
  signal rematch002_in_cmd_accm_inst_kernel_cmd_ready           : std_logic;
  signal rematch002_in_cmd_accm_inst_kernel_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch002_in_cmd_accm_inst_kernel_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch002_in_cmd_accm_inst_kernel_cmd_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch002_in_cmd_accm_inst_nucleus_cmd_valid          : std_logic;
  signal rematch002_in_cmd_accm_inst_nucleus_cmd_ready          : std_logic;
  signal rematch002_in_cmd_accm_inst_nucleus_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch002_in_cmd_accm_inst_nucleus_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch002_in_cmd_accm_inst_nucleus_cmd_ctrl           : std_logic_vector(2*REMATCH002_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch002_in_cmd_accm_inst_nucleus_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch003_in_cmd_accm_inst_kernel_cmd_valid           : std_logic;
  signal rematch003_in_cmd_accm_inst_kernel_cmd_ready           : std_logic;
  signal rematch003_in_cmd_accm_inst_kernel_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch003_in_cmd_accm_inst_kernel_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch003_in_cmd_accm_inst_kernel_cmd_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch003_in_cmd_accm_inst_nucleus_cmd_valid          : std_logic;
  signal rematch003_in_cmd_accm_inst_nucleus_cmd_ready          : std_logic;
  signal rematch003_in_cmd_accm_inst_nucleus_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch003_in_cmd_accm_inst_nucleus_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch003_in_cmd_accm_inst_nucleus_cmd_ctrl           : std_logic_vector(2*REMATCH003_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch003_in_cmd_accm_inst_nucleus_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch004_in_cmd_accm_inst_kernel_cmd_valid           : std_logic;
  signal rematch004_in_cmd_accm_inst_kernel_cmd_ready           : std_logic;
  signal rematch004_in_cmd_accm_inst_kernel_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch004_in_cmd_accm_inst_kernel_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch004_in_cmd_accm_inst_kernel_cmd_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch004_in_cmd_accm_inst_nucleus_cmd_valid          : std_logic;
  signal rematch004_in_cmd_accm_inst_nucleus_cmd_ready          : std_logic;
  signal rematch004_in_cmd_accm_inst_nucleus_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch004_in_cmd_accm_inst_nucleus_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch004_in_cmd_accm_inst_nucleus_cmd_ctrl           : std_logic_vector(2*REMATCH004_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch004_in_cmd_accm_inst_nucleus_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch005_in_cmd_accm_inst_kernel_cmd_valid           : std_logic;
  signal rematch005_in_cmd_accm_inst_kernel_cmd_ready           : std_logic;
  signal rematch005_in_cmd_accm_inst_kernel_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch005_in_cmd_accm_inst_kernel_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch005_in_cmd_accm_inst_kernel_cmd_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch005_in_cmd_accm_inst_nucleus_cmd_valid          : std_logic;
  signal rematch005_in_cmd_accm_inst_nucleus_cmd_ready          : std_logic;
  signal rematch005_in_cmd_accm_inst_nucleus_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch005_in_cmd_accm_inst_nucleus_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch005_in_cmd_accm_inst_nucleus_cmd_ctrl           : std_logic_vector(2*REMATCH005_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch005_in_cmd_accm_inst_nucleus_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch006_in_cmd_accm_inst_kernel_cmd_valid           : std_logic;
  signal rematch006_in_cmd_accm_inst_kernel_cmd_ready           : std_logic;
  signal rematch006_in_cmd_accm_inst_kernel_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch006_in_cmd_accm_inst_kernel_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch006_in_cmd_accm_inst_kernel_cmd_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch006_in_cmd_accm_inst_nucleus_cmd_valid          : std_logic;
  signal rematch006_in_cmd_accm_inst_nucleus_cmd_ready          : std_logic;
  signal rematch006_in_cmd_accm_inst_nucleus_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch006_in_cmd_accm_inst_nucleus_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch006_in_cmd_accm_inst_nucleus_cmd_ctrl           : std_logic_vector(2*REMATCH006_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch006_in_cmd_accm_inst_nucleus_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch007_in_cmd_accm_inst_kernel_cmd_valid           : std_logic;
  signal rematch007_in_cmd_accm_inst_kernel_cmd_ready           : std_logic;
  signal rematch007_in_cmd_accm_inst_kernel_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch007_in_cmd_accm_inst_kernel_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch007_in_cmd_accm_inst_kernel_cmd_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch007_in_cmd_accm_inst_nucleus_cmd_valid          : std_logic;
  signal rematch007_in_cmd_accm_inst_nucleus_cmd_ready          : std_logic;
  signal rematch007_in_cmd_accm_inst_nucleus_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch007_in_cmd_accm_inst_nucleus_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch007_in_cmd_accm_inst_nucleus_cmd_ctrl           : std_logic_vector(2*REMATCH007_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch007_in_cmd_accm_inst_nucleus_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch008_in_cmd_accm_inst_kernel_cmd_valid           : std_logic;
  signal rematch008_in_cmd_accm_inst_kernel_cmd_ready           : std_logic;
  signal rematch008_in_cmd_accm_inst_kernel_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch008_in_cmd_accm_inst_kernel_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch008_in_cmd_accm_inst_kernel_cmd_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch008_in_cmd_accm_inst_nucleus_cmd_valid          : std_logic;
  signal rematch008_in_cmd_accm_inst_nucleus_cmd_ready          : std_logic;
  signal rematch008_in_cmd_accm_inst_nucleus_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch008_in_cmd_accm_inst_nucleus_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch008_in_cmd_accm_inst_nucleus_cmd_ctrl           : std_logic_vector(2*REMATCH008_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch008_in_cmd_accm_inst_nucleus_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch009_in_cmd_accm_inst_kernel_cmd_valid           : std_logic;
  signal rematch009_in_cmd_accm_inst_kernel_cmd_ready           : std_logic;
  signal rematch009_in_cmd_accm_inst_kernel_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch009_in_cmd_accm_inst_kernel_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch009_in_cmd_accm_inst_kernel_cmd_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch009_in_cmd_accm_inst_nucleus_cmd_valid          : std_logic;
  signal rematch009_in_cmd_accm_inst_nucleus_cmd_ready          : std_logic;
  signal rematch009_in_cmd_accm_inst_nucleus_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch009_in_cmd_accm_inst_nucleus_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch009_in_cmd_accm_inst_nucleus_cmd_ctrl           : std_logic_vector(2*REMATCH009_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch009_in_cmd_accm_inst_nucleus_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch010_in_cmd_accm_inst_kernel_cmd_valid           : std_logic;
  signal rematch010_in_cmd_accm_inst_kernel_cmd_ready           : std_logic;
  signal rematch010_in_cmd_accm_inst_kernel_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch010_in_cmd_accm_inst_kernel_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch010_in_cmd_accm_inst_kernel_cmd_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch010_in_cmd_accm_inst_nucleus_cmd_valid          : std_logic;
  signal rematch010_in_cmd_accm_inst_nucleus_cmd_ready          : std_logic;
  signal rematch010_in_cmd_accm_inst_nucleus_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch010_in_cmd_accm_inst_nucleus_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch010_in_cmd_accm_inst_nucleus_cmd_ctrl           : std_logic_vector(2*REMATCH010_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch010_in_cmd_accm_inst_nucleus_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch011_in_cmd_accm_inst_kernel_cmd_valid           : std_logic;
  signal rematch011_in_cmd_accm_inst_kernel_cmd_ready           : std_logic;
  signal rematch011_in_cmd_accm_inst_kernel_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch011_in_cmd_accm_inst_kernel_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch011_in_cmd_accm_inst_kernel_cmd_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch011_in_cmd_accm_inst_nucleus_cmd_valid          : std_logic;
  signal rematch011_in_cmd_accm_inst_nucleus_cmd_ready          : std_logic;
  signal rematch011_in_cmd_accm_inst_nucleus_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch011_in_cmd_accm_inst_nucleus_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch011_in_cmd_accm_inst_nucleus_cmd_ctrl           : std_logic_vector(2*REMATCH011_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch011_in_cmd_accm_inst_nucleus_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch012_in_cmd_accm_inst_kernel_cmd_valid           : std_logic;
  signal rematch012_in_cmd_accm_inst_kernel_cmd_ready           : std_logic;
  signal rematch012_in_cmd_accm_inst_kernel_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch012_in_cmd_accm_inst_kernel_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch012_in_cmd_accm_inst_kernel_cmd_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch012_in_cmd_accm_inst_nucleus_cmd_valid          : std_logic;
  signal rematch012_in_cmd_accm_inst_nucleus_cmd_ready          : std_logic;
  signal rematch012_in_cmd_accm_inst_nucleus_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch012_in_cmd_accm_inst_nucleus_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch012_in_cmd_accm_inst_nucleus_cmd_ctrl           : std_logic_vector(2*REMATCH012_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch012_in_cmd_accm_inst_nucleus_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch013_in_cmd_accm_inst_kernel_cmd_valid           : std_logic;
  signal rematch013_in_cmd_accm_inst_kernel_cmd_ready           : std_logic;
  signal rematch013_in_cmd_accm_inst_kernel_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch013_in_cmd_accm_inst_kernel_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch013_in_cmd_accm_inst_kernel_cmd_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch013_in_cmd_accm_inst_nucleus_cmd_valid          : std_logic;
  signal rematch013_in_cmd_accm_inst_nucleus_cmd_ready          : std_logic;
  signal rematch013_in_cmd_accm_inst_nucleus_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch013_in_cmd_accm_inst_nucleus_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch013_in_cmd_accm_inst_nucleus_cmd_ctrl           : std_logic_vector(2*REMATCH013_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch013_in_cmd_accm_inst_nucleus_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch014_in_cmd_accm_inst_kernel_cmd_valid           : std_logic;
  signal rematch014_in_cmd_accm_inst_kernel_cmd_ready           : std_logic;
  signal rematch014_in_cmd_accm_inst_kernel_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch014_in_cmd_accm_inst_kernel_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch014_in_cmd_accm_inst_kernel_cmd_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch014_in_cmd_accm_inst_nucleus_cmd_valid          : std_logic;
  signal rematch014_in_cmd_accm_inst_nucleus_cmd_ready          : std_logic;
  signal rematch014_in_cmd_accm_inst_nucleus_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch014_in_cmd_accm_inst_nucleus_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch014_in_cmd_accm_inst_nucleus_cmd_ctrl           : std_logic_vector(2*REMATCH014_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch014_in_cmd_accm_inst_nucleus_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch015_in_cmd_accm_inst_kernel_cmd_valid           : std_logic;
  signal rematch015_in_cmd_accm_inst_kernel_cmd_ready           : std_logic;
  signal rematch015_in_cmd_accm_inst_kernel_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch015_in_cmd_accm_inst_kernel_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch015_in_cmd_accm_inst_kernel_cmd_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch015_in_cmd_accm_inst_nucleus_cmd_valid          : std_logic;
  signal rematch015_in_cmd_accm_inst_nucleus_cmd_ready          : std_logic;
  signal rematch015_in_cmd_accm_inst_nucleus_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch015_in_cmd_accm_inst_nucleus_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch015_in_cmd_accm_inst_nucleus_cmd_ctrl           : std_logic_vector(2*REMATCH015_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch015_in_cmd_accm_inst_nucleus_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch000_taxi_out_cmd_accm_inst_kernel_cmd_valid     : std_logic;
  signal rematch000_taxi_out_cmd_accm_inst_kernel_cmd_ready     : std_logic;
  signal rematch000_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch000_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch000_taxi_out_cmd_accm_inst_kernel_cmd_tag       : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch000_taxi_out_cmd_accm_inst_nucleus_cmd_valid    : std_logic;
  signal rematch000_taxi_out_cmd_accm_inst_nucleus_cmd_ready    : std_logic;
  signal rematch000_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch000_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch000_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl     : std_logic_vector(REMATCH000_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch000_taxi_out_cmd_accm_inst_nucleus_cmd_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch001_taxi_out_cmd_accm_inst_kernel_cmd_valid     : std_logic;
  signal rematch001_taxi_out_cmd_accm_inst_kernel_cmd_ready     : std_logic;
  signal rematch001_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch001_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch001_taxi_out_cmd_accm_inst_kernel_cmd_tag       : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch001_taxi_out_cmd_accm_inst_nucleus_cmd_valid    : std_logic;
  signal rematch001_taxi_out_cmd_accm_inst_nucleus_cmd_ready    : std_logic;
  signal rematch001_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch001_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch001_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl     : std_logic_vector(REMATCH001_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch001_taxi_out_cmd_accm_inst_nucleus_cmd_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch002_taxi_out_cmd_accm_inst_kernel_cmd_valid     : std_logic;
  signal rematch002_taxi_out_cmd_accm_inst_kernel_cmd_ready     : std_logic;
  signal rematch002_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch002_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch002_taxi_out_cmd_accm_inst_kernel_cmd_tag       : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch002_taxi_out_cmd_accm_inst_nucleus_cmd_valid    : std_logic;
  signal rematch002_taxi_out_cmd_accm_inst_nucleus_cmd_ready    : std_logic;
  signal rematch002_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch002_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch002_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl     : std_logic_vector(REMATCH002_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch002_taxi_out_cmd_accm_inst_nucleus_cmd_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch003_taxi_out_cmd_accm_inst_kernel_cmd_valid     : std_logic;
  signal rematch003_taxi_out_cmd_accm_inst_kernel_cmd_ready     : std_logic;
  signal rematch003_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch003_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch003_taxi_out_cmd_accm_inst_kernel_cmd_tag       : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch003_taxi_out_cmd_accm_inst_nucleus_cmd_valid    : std_logic;
  signal rematch003_taxi_out_cmd_accm_inst_nucleus_cmd_ready    : std_logic;
  signal rematch003_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch003_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch003_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl     : std_logic_vector(REMATCH003_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch003_taxi_out_cmd_accm_inst_nucleus_cmd_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch004_taxi_out_cmd_accm_inst_kernel_cmd_valid     : std_logic;
  signal rematch004_taxi_out_cmd_accm_inst_kernel_cmd_ready     : std_logic;
  signal rematch004_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch004_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch004_taxi_out_cmd_accm_inst_kernel_cmd_tag       : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch004_taxi_out_cmd_accm_inst_nucleus_cmd_valid    : std_logic;
  signal rematch004_taxi_out_cmd_accm_inst_nucleus_cmd_ready    : std_logic;
  signal rematch004_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch004_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch004_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl     : std_logic_vector(REMATCH004_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch004_taxi_out_cmd_accm_inst_nucleus_cmd_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch005_taxi_out_cmd_accm_inst_kernel_cmd_valid     : std_logic;
  signal rematch005_taxi_out_cmd_accm_inst_kernel_cmd_ready     : std_logic;
  signal rematch005_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch005_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch005_taxi_out_cmd_accm_inst_kernel_cmd_tag       : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch005_taxi_out_cmd_accm_inst_nucleus_cmd_valid    : std_logic;
  signal rematch005_taxi_out_cmd_accm_inst_nucleus_cmd_ready    : std_logic;
  signal rematch005_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch005_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch005_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl     : std_logic_vector(REMATCH005_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch005_taxi_out_cmd_accm_inst_nucleus_cmd_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch006_taxi_out_cmd_accm_inst_kernel_cmd_valid     : std_logic;
  signal rematch006_taxi_out_cmd_accm_inst_kernel_cmd_ready     : std_logic;
  signal rematch006_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch006_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch006_taxi_out_cmd_accm_inst_kernel_cmd_tag       : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch006_taxi_out_cmd_accm_inst_nucleus_cmd_valid    : std_logic;
  signal rematch006_taxi_out_cmd_accm_inst_nucleus_cmd_ready    : std_logic;
  signal rematch006_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch006_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch006_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl     : std_logic_vector(REMATCH006_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch006_taxi_out_cmd_accm_inst_nucleus_cmd_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch007_taxi_out_cmd_accm_inst_kernel_cmd_valid     : std_logic;
  signal rematch007_taxi_out_cmd_accm_inst_kernel_cmd_ready     : std_logic;
  signal rematch007_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch007_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch007_taxi_out_cmd_accm_inst_kernel_cmd_tag       : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch007_taxi_out_cmd_accm_inst_nucleus_cmd_valid    : std_logic;
  signal rematch007_taxi_out_cmd_accm_inst_nucleus_cmd_ready    : std_logic;
  signal rematch007_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch007_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch007_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl     : std_logic_vector(REMATCH007_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch007_taxi_out_cmd_accm_inst_nucleus_cmd_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch008_taxi_out_cmd_accm_inst_kernel_cmd_valid     : std_logic;
  signal rematch008_taxi_out_cmd_accm_inst_kernel_cmd_ready     : std_logic;
  signal rematch008_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch008_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch008_taxi_out_cmd_accm_inst_kernel_cmd_tag       : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch008_taxi_out_cmd_accm_inst_nucleus_cmd_valid    : std_logic;
  signal rematch008_taxi_out_cmd_accm_inst_nucleus_cmd_ready    : std_logic;
  signal rematch008_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch008_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch008_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl     : std_logic_vector(REMATCH008_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch008_taxi_out_cmd_accm_inst_nucleus_cmd_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch009_taxi_out_cmd_accm_inst_kernel_cmd_valid     : std_logic;
  signal rematch009_taxi_out_cmd_accm_inst_kernel_cmd_ready     : std_logic;
  signal rematch009_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch009_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch009_taxi_out_cmd_accm_inst_kernel_cmd_tag       : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch009_taxi_out_cmd_accm_inst_nucleus_cmd_valid    : std_logic;
  signal rematch009_taxi_out_cmd_accm_inst_nucleus_cmd_ready    : std_logic;
  signal rematch009_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch009_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch009_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl     : std_logic_vector(REMATCH009_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch009_taxi_out_cmd_accm_inst_nucleus_cmd_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch010_taxi_out_cmd_accm_inst_kernel_cmd_valid     : std_logic;
  signal rematch010_taxi_out_cmd_accm_inst_kernel_cmd_ready     : std_logic;
  signal rematch010_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch010_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch010_taxi_out_cmd_accm_inst_kernel_cmd_tag       : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch010_taxi_out_cmd_accm_inst_nucleus_cmd_valid    : std_logic;
  signal rematch010_taxi_out_cmd_accm_inst_nucleus_cmd_ready    : std_logic;
  signal rematch010_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch010_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch010_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl     : std_logic_vector(REMATCH010_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch010_taxi_out_cmd_accm_inst_nucleus_cmd_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch011_taxi_out_cmd_accm_inst_kernel_cmd_valid     : std_logic;
  signal rematch011_taxi_out_cmd_accm_inst_kernel_cmd_ready     : std_logic;
  signal rematch011_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch011_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch011_taxi_out_cmd_accm_inst_kernel_cmd_tag       : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch011_taxi_out_cmd_accm_inst_nucleus_cmd_valid    : std_logic;
  signal rematch011_taxi_out_cmd_accm_inst_nucleus_cmd_ready    : std_logic;
  signal rematch011_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch011_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch011_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl     : std_logic_vector(REMATCH011_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch011_taxi_out_cmd_accm_inst_nucleus_cmd_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch012_taxi_out_cmd_accm_inst_kernel_cmd_valid     : std_logic;
  signal rematch012_taxi_out_cmd_accm_inst_kernel_cmd_ready     : std_logic;
  signal rematch012_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch012_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch012_taxi_out_cmd_accm_inst_kernel_cmd_tag       : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch012_taxi_out_cmd_accm_inst_nucleus_cmd_valid    : std_logic;
  signal rematch012_taxi_out_cmd_accm_inst_nucleus_cmd_ready    : std_logic;
  signal rematch012_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch012_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch012_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl     : std_logic_vector(REMATCH012_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch012_taxi_out_cmd_accm_inst_nucleus_cmd_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch013_taxi_out_cmd_accm_inst_kernel_cmd_valid     : std_logic;
  signal rematch013_taxi_out_cmd_accm_inst_kernel_cmd_ready     : std_logic;
  signal rematch013_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch013_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch013_taxi_out_cmd_accm_inst_kernel_cmd_tag       : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch013_taxi_out_cmd_accm_inst_nucleus_cmd_valid    : std_logic;
  signal rematch013_taxi_out_cmd_accm_inst_nucleus_cmd_ready    : std_logic;
  signal rematch013_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch013_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch013_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl     : std_logic_vector(REMATCH013_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch013_taxi_out_cmd_accm_inst_nucleus_cmd_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch014_taxi_out_cmd_accm_inst_kernel_cmd_valid     : std_logic;
  signal rematch014_taxi_out_cmd_accm_inst_kernel_cmd_ready     : std_logic;
  signal rematch014_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch014_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch014_taxi_out_cmd_accm_inst_kernel_cmd_tag       : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch014_taxi_out_cmd_accm_inst_nucleus_cmd_valid    : std_logic;
  signal rematch014_taxi_out_cmd_accm_inst_nucleus_cmd_ready    : std_logic;
  signal rematch014_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch014_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch014_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl     : std_logic_vector(REMATCH014_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch014_taxi_out_cmd_accm_inst_nucleus_cmd_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch015_taxi_out_cmd_accm_inst_kernel_cmd_valid     : std_logic;
  signal rematch015_taxi_out_cmd_accm_inst_kernel_cmd_ready     : std_logic;
  signal rematch015_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch015_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch015_taxi_out_cmd_accm_inst_kernel_cmd_tag       : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch015_taxi_out_cmd_accm_inst_nucleus_cmd_valid    : std_logic;
  signal rematch015_taxi_out_cmd_accm_inst_nucleus_cmd_ready    : std_logic;
  signal rematch015_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch015_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal rematch015_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl     : std_logic_vector(REMATCH015_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch015_taxi_out_cmd_accm_inst_nucleus_cmd_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal rematch000_in_cmd_accm_inst_ctrl       : std_logic_vector(2*REMATCH000_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch001_in_cmd_accm_inst_ctrl       : std_logic_vector(2*REMATCH001_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch002_in_cmd_accm_inst_ctrl       : std_logic_vector(2*REMATCH002_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch003_in_cmd_accm_inst_ctrl       : std_logic_vector(2*REMATCH003_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch004_in_cmd_accm_inst_ctrl       : std_logic_vector(2*REMATCH004_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch005_in_cmd_accm_inst_ctrl       : std_logic_vector(2*REMATCH005_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch006_in_cmd_accm_inst_ctrl       : std_logic_vector(2*REMATCH006_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch007_in_cmd_accm_inst_ctrl       : std_logic_vector(2*REMATCH007_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch008_in_cmd_accm_inst_ctrl       : std_logic_vector(2*REMATCH008_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch009_in_cmd_accm_inst_ctrl       : std_logic_vector(2*REMATCH009_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch010_in_cmd_accm_inst_ctrl       : std_logic_vector(2*REMATCH010_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch011_in_cmd_accm_inst_ctrl       : std_logic_vector(2*REMATCH011_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch012_in_cmd_accm_inst_ctrl       : std_logic_vector(2*REMATCH012_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch013_in_cmd_accm_inst_ctrl       : std_logic_vector(2*REMATCH013_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch014_in_cmd_accm_inst_ctrl       : std_logic_vector(2*REMATCH014_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch015_in_cmd_accm_inst_ctrl       : std_logic_vector(2*REMATCH015_IN_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch000_taxi_out_cmd_accm_inst_ctrl : std_logic_vector(REMATCH000_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch001_taxi_out_cmd_accm_inst_ctrl : std_logic_vector(REMATCH001_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch002_taxi_out_cmd_accm_inst_ctrl : std_logic_vector(REMATCH002_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch003_taxi_out_cmd_accm_inst_ctrl : std_logic_vector(REMATCH003_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch004_taxi_out_cmd_accm_inst_ctrl : std_logic_vector(REMATCH004_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch005_taxi_out_cmd_accm_inst_ctrl : std_logic_vector(REMATCH005_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch006_taxi_out_cmd_accm_inst_ctrl : std_logic_vector(REMATCH006_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch007_taxi_out_cmd_accm_inst_ctrl : std_logic_vector(REMATCH007_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch008_taxi_out_cmd_accm_inst_ctrl : std_logic_vector(REMATCH008_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch009_taxi_out_cmd_accm_inst_ctrl : std_logic_vector(REMATCH009_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch010_taxi_out_cmd_accm_inst_ctrl : std_logic_vector(REMATCH010_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch011_taxi_out_cmd_accm_inst_ctrl : std_logic_vector(REMATCH011_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch012_taxi_out_cmd_accm_inst_ctrl : std_logic_vector(REMATCH012_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch013_taxi_out_cmd_accm_inst_ctrl : std_logic_vector(REMATCH013_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch014_taxi_out_cmd_accm_inst_ctrl : std_logic_vector(REMATCH014_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);
  signal rematch015_taxi_out_cmd_accm_inst_ctrl : std_logic_vector(REMATCH015_TAXI_OUT_BUS_ADDR_WIDTH-1 downto 0);

begin
  Kernel_inst : Kernel
    generic map (
      INDEX_WIDTH => 32,
      TAG_WIDTH   => 1
    )
    port map (
      kcd_clk                          => kcd_clk,
      kcd_reset                        => kcd_reset,
      rematch000_in_valid              => Kernel_inst_rematch000_in_valid,
      rematch000_in_ready              => Kernel_inst_rematch000_in_ready,
      rematch000_in_dvalid             => Kernel_inst_rematch000_in_dvalid,
      rematch000_in_last               => Kernel_inst_rematch000_in_last,
      rematch000_in_length             => Kernel_inst_rematch000_in_length,
      rematch000_in_count              => Kernel_inst_rematch000_in_count,
      rematch000_in_chars_valid        => Kernel_inst_rematch000_in_chars_valid,
      rematch000_in_chars_ready        => Kernel_inst_rematch000_in_chars_ready,
      rematch000_in_chars_dvalid       => Kernel_inst_rematch000_in_chars_dvalid,
      rematch000_in_chars_last         => Kernel_inst_rematch000_in_chars_last,
      rematch000_in_chars              => Kernel_inst_rematch000_in_chars,
      rematch000_in_chars_count        => Kernel_inst_rematch000_in_chars_count,
      rematch000_in_unl_valid          => Kernel_inst_rematch000_in_unl_valid,
      rematch000_in_unl_ready          => Kernel_inst_rematch000_in_unl_ready,
      rematch000_in_unl_tag            => Kernel_inst_rematch000_in_unl_tag,
      rematch000_in_cmd_valid          => Kernel_inst_rematch000_in_cmd_valid,
      rematch000_in_cmd_ready          => Kernel_inst_rematch000_in_cmd_ready,
      rematch000_in_cmd_firstIdx       => Kernel_inst_rematch000_in_cmd_firstIdx,
      rematch000_in_cmd_lastIdx        => Kernel_inst_rematch000_in_cmd_lastIdx,
      rematch000_in_cmd_tag            => Kernel_inst_rematch000_in_cmd_tag,
      rematch001_in_valid              => Kernel_inst_rematch001_in_valid,
      rematch001_in_ready              => Kernel_inst_rematch001_in_ready,
      rematch001_in_dvalid             => Kernel_inst_rematch001_in_dvalid,
      rematch001_in_last               => Kernel_inst_rematch001_in_last,
      rematch001_in_length             => Kernel_inst_rematch001_in_length,
      rematch001_in_count              => Kernel_inst_rematch001_in_count,
      rematch001_in_chars_valid        => Kernel_inst_rematch001_in_chars_valid,
      rematch001_in_chars_ready        => Kernel_inst_rematch001_in_chars_ready,
      rematch001_in_chars_dvalid       => Kernel_inst_rematch001_in_chars_dvalid,
      rematch001_in_chars_last         => Kernel_inst_rematch001_in_chars_last,
      rematch001_in_chars              => Kernel_inst_rematch001_in_chars,
      rematch001_in_chars_count        => Kernel_inst_rematch001_in_chars_count,
      rematch001_in_unl_valid          => Kernel_inst_rematch001_in_unl_valid,
      rematch001_in_unl_ready          => Kernel_inst_rematch001_in_unl_ready,
      rematch001_in_unl_tag            => Kernel_inst_rematch001_in_unl_tag,
      rematch001_in_cmd_valid          => Kernel_inst_rematch001_in_cmd_valid,
      rematch001_in_cmd_ready          => Kernel_inst_rematch001_in_cmd_ready,
      rematch001_in_cmd_firstIdx       => Kernel_inst_rematch001_in_cmd_firstIdx,
      rematch001_in_cmd_lastIdx        => Kernel_inst_rematch001_in_cmd_lastIdx,
      rematch001_in_cmd_tag            => Kernel_inst_rematch001_in_cmd_tag,
      rematch002_in_valid              => Kernel_inst_rematch002_in_valid,
      rematch002_in_ready              => Kernel_inst_rematch002_in_ready,
      rematch002_in_dvalid             => Kernel_inst_rematch002_in_dvalid,
      rematch002_in_last               => Kernel_inst_rematch002_in_last,
      rematch002_in_length             => Kernel_inst_rematch002_in_length,
      rematch002_in_count              => Kernel_inst_rematch002_in_count,
      rematch002_in_chars_valid        => Kernel_inst_rematch002_in_chars_valid,
      rematch002_in_chars_ready        => Kernel_inst_rematch002_in_chars_ready,
      rematch002_in_chars_dvalid       => Kernel_inst_rematch002_in_chars_dvalid,
      rematch002_in_chars_last         => Kernel_inst_rematch002_in_chars_last,
      rematch002_in_chars              => Kernel_inst_rematch002_in_chars,
      rematch002_in_chars_count        => Kernel_inst_rematch002_in_chars_count,
      rematch002_in_unl_valid          => Kernel_inst_rematch002_in_unl_valid,
      rematch002_in_unl_ready          => Kernel_inst_rematch002_in_unl_ready,
      rematch002_in_unl_tag            => Kernel_inst_rematch002_in_unl_tag,
      rematch002_in_cmd_valid          => Kernel_inst_rematch002_in_cmd_valid,
      rematch002_in_cmd_ready          => Kernel_inst_rematch002_in_cmd_ready,
      rematch002_in_cmd_firstIdx       => Kernel_inst_rematch002_in_cmd_firstIdx,
      rematch002_in_cmd_lastIdx        => Kernel_inst_rematch002_in_cmd_lastIdx,
      rematch002_in_cmd_tag            => Kernel_inst_rematch002_in_cmd_tag,
      rematch003_in_valid              => Kernel_inst_rematch003_in_valid,
      rematch003_in_ready              => Kernel_inst_rematch003_in_ready,
      rematch003_in_dvalid             => Kernel_inst_rematch003_in_dvalid,
      rematch003_in_last               => Kernel_inst_rematch003_in_last,
      rematch003_in_length             => Kernel_inst_rematch003_in_length,
      rematch003_in_count              => Kernel_inst_rematch003_in_count,
      rematch003_in_chars_valid        => Kernel_inst_rematch003_in_chars_valid,
      rematch003_in_chars_ready        => Kernel_inst_rematch003_in_chars_ready,
      rematch003_in_chars_dvalid       => Kernel_inst_rematch003_in_chars_dvalid,
      rematch003_in_chars_last         => Kernel_inst_rematch003_in_chars_last,
      rematch003_in_chars              => Kernel_inst_rematch003_in_chars,
      rematch003_in_chars_count        => Kernel_inst_rematch003_in_chars_count,
      rematch003_in_unl_valid          => Kernel_inst_rematch003_in_unl_valid,
      rematch003_in_unl_ready          => Kernel_inst_rematch003_in_unl_ready,
      rematch003_in_unl_tag            => Kernel_inst_rematch003_in_unl_tag,
      rematch003_in_cmd_valid          => Kernel_inst_rematch003_in_cmd_valid,
      rematch003_in_cmd_ready          => Kernel_inst_rematch003_in_cmd_ready,
      rematch003_in_cmd_firstIdx       => Kernel_inst_rematch003_in_cmd_firstIdx,
      rematch003_in_cmd_lastIdx        => Kernel_inst_rematch003_in_cmd_lastIdx,
      rematch003_in_cmd_tag            => Kernel_inst_rematch003_in_cmd_tag,
      rematch004_in_valid              => Kernel_inst_rematch004_in_valid,
      rematch004_in_ready              => Kernel_inst_rematch004_in_ready,
      rematch004_in_dvalid             => Kernel_inst_rematch004_in_dvalid,
      rematch004_in_last               => Kernel_inst_rematch004_in_last,
      rematch004_in_length             => Kernel_inst_rematch004_in_length,
      rematch004_in_count              => Kernel_inst_rematch004_in_count,
      rematch004_in_chars_valid        => Kernel_inst_rematch004_in_chars_valid,
      rematch004_in_chars_ready        => Kernel_inst_rematch004_in_chars_ready,
      rematch004_in_chars_dvalid       => Kernel_inst_rematch004_in_chars_dvalid,
      rematch004_in_chars_last         => Kernel_inst_rematch004_in_chars_last,
      rematch004_in_chars              => Kernel_inst_rematch004_in_chars,
      rematch004_in_chars_count        => Kernel_inst_rematch004_in_chars_count,
      rematch004_in_unl_valid          => Kernel_inst_rematch004_in_unl_valid,
      rematch004_in_unl_ready          => Kernel_inst_rematch004_in_unl_ready,
      rematch004_in_unl_tag            => Kernel_inst_rematch004_in_unl_tag,
      rematch004_in_cmd_valid          => Kernel_inst_rematch004_in_cmd_valid,
      rematch004_in_cmd_ready          => Kernel_inst_rematch004_in_cmd_ready,
      rematch004_in_cmd_firstIdx       => Kernel_inst_rematch004_in_cmd_firstIdx,
      rematch004_in_cmd_lastIdx        => Kernel_inst_rematch004_in_cmd_lastIdx,
      rematch004_in_cmd_tag            => Kernel_inst_rematch004_in_cmd_tag,
      rematch005_in_valid              => Kernel_inst_rematch005_in_valid,
      rematch005_in_ready              => Kernel_inst_rematch005_in_ready,
      rematch005_in_dvalid             => Kernel_inst_rematch005_in_dvalid,
      rematch005_in_last               => Kernel_inst_rematch005_in_last,
      rematch005_in_length             => Kernel_inst_rematch005_in_length,
      rematch005_in_count              => Kernel_inst_rematch005_in_count,
      rematch005_in_chars_valid        => Kernel_inst_rematch005_in_chars_valid,
      rematch005_in_chars_ready        => Kernel_inst_rematch005_in_chars_ready,
      rematch005_in_chars_dvalid       => Kernel_inst_rematch005_in_chars_dvalid,
      rematch005_in_chars_last         => Kernel_inst_rematch005_in_chars_last,
      rematch005_in_chars              => Kernel_inst_rematch005_in_chars,
      rematch005_in_chars_count        => Kernel_inst_rematch005_in_chars_count,
      rematch005_in_unl_valid          => Kernel_inst_rematch005_in_unl_valid,
      rematch005_in_unl_ready          => Kernel_inst_rematch005_in_unl_ready,
      rematch005_in_unl_tag            => Kernel_inst_rematch005_in_unl_tag,
      rematch005_in_cmd_valid          => Kernel_inst_rematch005_in_cmd_valid,
      rematch005_in_cmd_ready          => Kernel_inst_rematch005_in_cmd_ready,
      rematch005_in_cmd_firstIdx       => Kernel_inst_rematch005_in_cmd_firstIdx,
      rematch005_in_cmd_lastIdx        => Kernel_inst_rematch005_in_cmd_lastIdx,
      rematch005_in_cmd_tag            => Kernel_inst_rematch005_in_cmd_tag,
      rematch006_in_valid              => Kernel_inst_rematch006_in_valid,
      rematch006_in_ready              => Kernel_inst_rematch006_in_ready,
      rematch006_in_dvalid             => Kernel_inst_rematch006_in_dvalid,
      rematch006_in_last               => Kernel_inst_rematch006_in_last,
      rematch006_in_length             => Kernel_inst_rematch006_in_length,
      rematch006_in_count              => Kernel_inst_rematch006_in_count,
      rematch006_in_chars_valid        => Kernel_inst_rematch006_in_chars_valid,
      rematch006_in_chars_ready        => Kernel_inst_rematch006_in_chars_ready,
      rematch006_in_chars_dvalid       => Kernel_inst_rematch006_in_chars_dvalid,
      rematch006_in_chars_last         => Kernel_inst_rematch006_in_chars_last,
      rematch006_in_chars              => Kernel_inst_rematch006_in_chars,
      rematch006_in_chars_count        => Kernel_inst_rematch006_in_chars_count,
      rematch006_in_unl_valid          => Kernel_inst_rematch006_in_unl_valid,
      rematch006_in_unl_ready          => Kernel_inst_rematch006_in_unl_ready,
      rematch006_in_unl_tag            => Kernel_inst_rematch006_in_unl_tag,
      rematch006_in_cmd_valid          => Kernel_inst_rematch006_in_cmd_valid,
      rematch006_in_cmd_ready          => Kernel_inst_rematch006_in_cmd_ready,
      rematch006_in_cmd_firstIdx       => Kernel_inst_rematch006_in_cmd_firstIdx,
      rematch006_in_cmd_lastIdx        => Kernel_inst_rematch006_in_cmd_lastIdx,
      rematch006_in_cmd_tag            => Kernel_inst_rematch006_in_cmd_tag,
      rematch007_in_valid              => Kernel_inst_rematch007_in_valid,
      rematch007_in_ready              => Kernel_inst_rematch007_in_ready,
      rematch007_in_dvalid             => Kernel_inst_rematch007_in_dvalid,
      rematch007_in_last               => Kernel_inst_rematch007_in_last,
      rematch007_in_length             => Kernel_inst_rematch007_in_length,
      rematch007_in_count              => Kernel_inst_rematch007_in_count,
      rematch007_in_chars_valid        => Kernel_inst_rematch007_in_chars_valid,
      rematch007_in_chars_ready        => Kernel_inst_rematch007_in_chars_ready,
      rematch007_in_chars_dvalid       => Kernel_inst_rematch007_in_chars_dvalid,
      rematch007_in_chars_last         => Kernel_inst_rematch007_in_chars_last,
      rematch007_in_chars              => Kernel_inst_rematch007_in_chars,
      rematch007_in_chars_count        => Kernel_inst_rematch007_in_chars_count,
      rematch007_in_unl_valid          => Kernel_inst_rematch007_in_unl_valid,
      rematch007_in_unl_ready          => Kernel_inst_rematch007_in_unl_ready,
      rematch007_in_unl_tag            => Kernel_inst_rematch007_in_unl_tag,
      rematch007_in_cmd_valid          => Kernel_inst_rematch007_in_cmd_valid,
      rematch007_in_cmd_ready          => Kernel_inst_rematch007_in_cmd_ready,
      rematch007_in_cmd_firstIdx       => Kernel_inst_rematch007_in_cmd_firstIdx,
      rematch007_in_cmd_lastIdx        => Kernel_inst_rematch007_in_cmd_lastIdx,
      rematch007_in_cmd_tag            => Kernel_inst_rematch007_in_cmd_tag,
      rematch008_in_valid              => Kernel_inst_rematch008_in_valid,
      rematch008_in_ready              => Kernel_inst_rematch008_in_ready,
      rematch008_in_dvalid             => Kernel_inst_rematch008_in_dvalid,
      rematch008_in_last               => Kernel_inst_rematch008_in_last,
      rematch008_in_length             => Kernel_inst_rematch008_in_length,
      rematch008_in_count              => Kernel_inst_rematch008_in_count,
      rematch008_in_chars_valid        => Kernel_inst_rematch008_in_chars_valid,
      rematch008_in_chars_ready        => Kernel_inst_rematch008_in_chars_ready,
      rematch008_in_chars_dvalid       => Kernel_inst_rematch008_in_chars_dvalid,
      rematch008_in_chars_last         => Kernel_inst_rematch008_in_chars_last,
      rematch008_in_chars              => Kernel_inst_rematch008_in_chars,
      rematch008_in_chars_count        => Kernel_inst_rematch008_in_chars_count,
      rematch008_in_unl_valid          => Kernel_inst_rematch008_in_unl_valid,
      rematch008_in_unl_ready          => Kernel_inst_rematch008_in_unl_ready,
      rematch008_in_unl_tag            => Kernel_inst_rematch008_in_unl_tag,
      rematch008_in_cmd_valid          => Kernel_inst_rematch008_in_cmd_valid,
      rematch008_in_cmd_ready          => Kernel_inst_rematch008_in_cmd_ready,
      rematch008_in_cmd_firstIdx       => Kernel_inst_rematch008_in_cmd_firstIdx,
      rematch008_in_cmd_lastIdx        => Kernel_inst_rematch008_in_cmd_lastIdx,
      rematch008_in_cmd_tag            => Kernel_inst_rematch008_in_cmd_tag,
      rematch009_in_valid              => Kernel_inst_rematch009_in_valid,
      rematch009_in_ready              => Kernel_inst_rematch009_in_ready,
      rematch009_in_dvalid             => Kernel_inst_rematch009_in_dvalid,
      rematch009_in_last               => Kernel_inst_rematch009_in_last,
      rematch009_in_length             => Kernel_inst_rematch009_in_length,
      rematch009_in_count              => Kernel_inst_rematch009_in_count,
      rematch009_in_chars_valid        => Kernel_inst_rematch009_in_chars_valid,
      rematch009_in_chars_ready        => Kernel_inst_rematch009_in_chars_ready,
      rematch009_in_chars_dvalid       => Kernel_inst_rematch009_in_chars_dvalid,
      rematch009_in_chars_last         => Kernel_inst_rematch009_in_chars_last,
      rematch009_in_chars              => Kernel_inst_rematch009_in_chars,
      rematch009_in_chars_count        => Kernel_inst_rematch009_in_chars_count,
      rematch009_in_unl_valid          => Kernel_inst_rematch009_in_unl_valid,
      rematch009_in_unl_ready          => Kernel_inst_rematch009_in_unl_ready,
      rematch009_in_unl_tag            => Kernel_inst_rematch009_in_unl_tag,
      rematch009_in_cmd_valid          => Kernel_inst_rematch009_in_cmd_valid,
      rematch009_in_cmd_ready          => Kernel_inst_rematch009_in_cmd_ready,
      rematch009_in_cmd_firstIdx       => Kernel_inst_rematch009_in_cmd_firstIdx,
      rematch009_in_cmd_lastIdx        => Kernel_inst_rematch009_in_cmd_lastIdx,
      rematch009_in_cmd_tag            => Kernel_inst_rematch009_in_cmd_tag,
      rematch010_in_valid              => Kernel_inst_rematch010_in_valid,
      rematch010_in_ready              => Kernel_inst_rematch010_in_ready,
      rematch010_in_dvalid             => Kernel_inst_rematch010_in_dvalid,
      rematch010_in_last               => Kernel_inst_rematch010_in_last,
      rematch010_in_length             => Kernel_inst_rematch010_in_length,
      rematch010_in_count              => Kernel_inst_rematch010_in_count,
      rematch010_in_chars_valid        => Kernel_inst_rematch010_in_chars_valid,
      rematch010_in_chars_ready        => Kernel_inst_rematch010_in_chars_ready,
      rematch010_in_chars_dvalid       => Kernel_inst_rematch010_in_chars_dvalid,
      rematch010_in_chars_last         => Kernel_inst_rematch010_in_chars_last,
      rematch010_in_chars              => Kernel_inst_rematch010_in_chars,
      rematch010_in_chars_count        => Kernel_inst_rematch010_in_chars_count,
      rematch010_in_unl_valid          => Kernel_inst_rematch010_in_unl_valid,
      rematch010_in_unl_ready          => Kernel_inst_rematch010_in_unl_ready,
      rematch010_in_unl_tag            => Kernel_inst_rematch010_in_unl_tag,
      rematch010_in_cmd_valid          => Kernel_inst_rematch010_in_cmd_valid,
      rematch010_in_cmd_ready          => Kernel_inst_rematch010_in_cmd_ready,
      rematch010_in_cmd_firstIdx       => Kernel_inst_rematch010_in_cmd_firstIdx,
      rematch010_in_cmd_lastIdx        => Kernel_inst_rematch010_in_cmd_lastIdx,
      rematch010_in_cmd_tag            => Kernel_inst_rematch010_in_cmd_tag,
      rematch011_in_valid              => Kernel_inst_rematch011_in_valid,
      rematch011_in_ready              => Kernel_inst_rematch011_in_ready,
      rematch011_in_dvalid             => Kernel_inst_rematch011_in_dvalid,
      rematch011_in_last               => Kernel_inst_rematch011_in_last,
      rematch011_in_length             => Kernel_inst_rematch011_in_length,
      rematch011_in_count              => Kernel_inst_rematch011_in_count,
      rematch011_in_chars_valid        => Kernel_inst_rematch011_in_chars_valid,
      rematch011_in_chars_ready        => Kernel_inst_rematch011_in_chars_ready,
      rematch011_in_chars_dvalid       => Kernel_inst_rematch011_in_chars_dvalid,
      rematch011_in_chars_last         => Kernel_inst_rematch011_in_chars_last,
      rematch011_in_chars              => Kernel_inst_rematch011_in_chars,
      rematch011_in_chars_count        => Kernel_inst_rematch011_in_chars_count,
      rematch011_in_unl_valid          => Kernel_inst_rematch011_in_unl_valid,
      rematch011_in_unl_ready          => Kernel_inst_rematch011_in_unl_ready,
      rematch011_in_unl_tag            => Kernel_inst_rematch011_in_unl_tag,
      rematch011_in_cmd_valid          => Kernel_inst_rematch011_in_cmd_valid,
      rematch011_in_cmd_ready          => Kernel_inst_rematch011_in_cmd_ready,
      rematch011_in_cmd_firstIdx       => Kernel_inst_rematch011_in_cmd_firstIdx,
      rematch011_in_cmd_lastIdx        => Kernel_inst_rematch011_in_cmd_lastIdx,
      rematch011_in_cmd_tag            => Kernel_inst_rematch011_in_cmd_tag,
      rematch012_in_valid              => Kernel_inst_rematch012_in_valid,
      rematch012_in_ready              => Kernel_inst_rematch012_in_ready,
      rematch012_in_dvalid             => Kernel_inst_rematch012_in_dvalid,
      rematch012_in_last               => Kernel_inst_rematch012_in_last,
      rematch012_in_length             => Kernel_inst_rematch012_in_length,
      rematch012_in_count              => Kernel_inst_rematch012_in_count,
      rematch012_in_chars_valid        => Kernel_inst_rematch012_in_chars_valid,
      rematch012_in_chars_ready        => Kernel_inst_rematch012_in_chars_ready,
      rematch012_in_chars_dvalid       => Kernel_inst_rematch012_in_chars_dvalid,
      rematch012_in_chars_last         => Kernel_inst_rematch012_in_chars_last,
      rematch012_in_chars              => Kernel_inst_rematch012_in_chars,
      rematch012_in_chars_count        => Kernel_inst_rematch012_in_chars_count,
      rematch012_in_unl_valid          => Kernel_inst_rematch012_in_unl_valid,
      rematch012_in_unl_ready          => Kernel_inst_rematch012_in_unl_ready,
      rematch012_in_unl_tag            => Kernel_inst_rematch012_in_unl_tag,
      rematch012_in_cmd_valid          => Kernel_inst_rematch012_in_cmd_valid,
      rematch012_in_cmd_ready          => Kernel_inst_rematch012_in_cmd_ready,
      rematch012_in_cmd_firstIdx       => Kernel_inst_rematch012_in_cmd_firstIdx,
      rematch012_in_cmd_lastIdx        => Kernel_inst_rematch012_in_cmd_lastIdx,
      rematch012_in_cmd_tag            => Kernel_inst_rematch012_in_cmd_tag,
      rematch013_in_valid              => Kernel_inst_rematch013_in_valid,
      rematch013_in_ready              => Kernel_inst_rematch013_in_ready,
      rematch013_in_dvalid             => Kernel_inst_rematch013_in_dvalid,
      rematch013_in_last               => Kernel_inst_rematch013_in_last,
      rematch013_in_length             => Kernel_inst_rematch013_in_length,
      rematch013_in_count              => Kernel_inst_rematch013_in_count,
      rematch013_in_chars_valid        => Kernel_inst_rematch013_in_chars_valid,
      rematch013_in_chars_ready        => Kernel_inst_rematch013_in_chars_ready,
      rematch013_in_chars_dvalid       => Kernel_inst_rematch013_in_chars_dvalid,
      rematch013_in_chars_last         => Kernel_inst_rematch013_in_chars_last,
      rematch013_in_chars              => Kernel_inst_rematch013_in_chars,
      rematch013_in_chars_count        => Kernel_inst_rematch013_in_chars_count,
      rematch013_in_unl_valid          => Kernel_inst_rematch013_in_unl_valid,
      rematch013_in_unl_ready          => Kernel_inst_rematch013_in_unl_ready,
      rematch013_in_unl_tag            => Kernel_inst_rematch013_in_unl_tag,
      rematch013_in_cmd_valid          => Kernel_inst_rematch013_in_cmd_valid,
      rematch013_in_cmd_ready          => Kernel_inst_rematch013_in_cmd_ready,
      rematch013_in_cmd_firstIdx       => Kernel_inst_rematch013_in_cmd_firstIdx,
      rematch013_in_cmd_lastIdx        => Kernel_inst_rematch013_in_cmd_lastIdx,
      rematch013_in_cmd_tag            => Kernel_inst_rematch013_in_cmd_tag,
      rematch014_in_valid              => Kernel_inst_rematch014_in_valid,
      rematch014_in_ready              => Kernel_inst_rematch014_in_ready,
      rematch014_in_dvalid             => Kernel_inst_rematch014_in_dvalid,
      rematch014_in_last               => Kernel_inst_rematch014_in_last,
      rematch014_in_length             => Kernel_inst_rematch014_in_length,
      rematch014_in_count              => Kernel_inst_rematch014_in_count,
      rematch014_in_chars_valid        => Kernel_inst_rematch014_in_chars_valid,
      rematch014_in_chars_ready        => Kernel_inst_rematch014_in_chars_ready,
      rematch014_in_chars_dvalid       => Kernel_inst_rematch014_in_chars_dvalid,
      rematch014_in_chars_last         => Kernel_inst_rematch014_in_chars_last,
      rematch014_in_chars              => Kernel_inst_rematch014_in_chars,
      rematch014_in_chars_count        => Kernel_inst_rematch014_in_chars_count,
      rematch014_in_unl_valid          => Kernel_inst_rematch014_in_unl_valid,
      rematch014_in_unl_ready          => Kernel_inst_rematch014_in_unl_ready,
      rematch014_in_unl_tag            => Kernel_inst_rematch014_in_unl_tag,
      rematch014_in_cmd_valid          => Kernel_inst_rematch014_in_cmd_valid,
      rematch014_in_cmd_ready          => Kernel_inst_rematch014_in_cmd_ready,
      rematch014_in_cmd_firstIdx       => Kernel_inst_rematch014_in_cmd_firstIdx,
      rematch014_in_cmd_lastIdx        => Kernel_inst_rematch014_in_cmd_lastIdx,
      rematch014_in_cmd_tag            => Kernel_inst_rematch014_in_cmd_tag,
      rematch015_in_valid              => Kernel_inst_rematch015_in_valid,
      rematch015_in_ready              => Kernel_inst_rematch015_in_ready,
      rematch015_in_dvalid             => Kernel_inst_rematch015_in_dvalid,
      rematch015_in_last               => Kernel_inst_rematch015_in_last,
      rematch015_in_length             => Kernel_inst_rematch015_in_length,
      rematch015_in_count              => Kernel_inst_rematch015_in_count,
      rematch015_in_chars_valid        => Kernel_inst_rematch015_in_chars_valid,
      rematch015_in_chars_ready        => Kernel_inst_rematch015_in_chars_ready,
      rematch015_in_chars_dvalid       => Kernel_inst_rematch015_in_chars_dvalid,
      rematch015_in_chars_last         => Kernel_inst_rematch015_in_chars_last,
      rematch015_in_chars              => Kernel_inst_rematch015_in_chars,
      rematch015_in_chars_count        => Kernel_inst_rematch015_in_chars_count,
      rematch015_in_unl_valid          => Kernel_inst_rematch015_in_unl_valid,
      rematch015_in_unl_ready          => Kernel_inst_rematch015_in_unl_ready,
      rematch015_in_unl_tag            => Kernel_inst_rematch015_in_unl_tag,
      rematch015_in_cmd_valid          => Kernel_inst_rematch015_in_cmd_valid,
      rematch015_in_cmd_ready          => Kernel_inst_rematch015_in_cmd_ready,
      rematch015_in_cmd_firstIdx       => Kernel_inst_rematch015_in_cmd_firstIdx,
      rematch015_in_cmd_lastIdx        => Kernel_inst_rematch015_in_cmd_lastIdx,
      rematch015_in_cmd_tag            => Kernel_inst_rematch015_in_cmd_tag,
      rematch000_taxi_out_valid        => Kernel_inst_rematch000_taxi_out_valid,
      rematch000_taxi_out_ready        => Kernel_inst_rematch000_taxi_out_ready,
      rematch000_taxi_out_dvalid       => Kernel_inst_rematch000_taxi_out_dvalid,
      rematch000_taxi_out_last         => Kernel_inst_rematch000_taxi_out_last,
      rematch000_taxi_out              => Kernel_inst_rematch000_taxi_out,
      rematch000_taxi_out_unl_valid    => Kernel_inst_rematch000_taxi_out_unl_valid,
      rematch000_taxi_out_unl_ready    => Kernel_inst_rematch000_taxi_out_unl_ready,
      rematch000_taxi_out_unl_tag      => Kernel_inst_rematch000_taxi_out_unl_tag,
      rematch000_taxi_out_cmd_valid    => Kernel_inst_rematch000_taxi_out_cmd_valid,
      rematch000_taxi_out_cmd_ready    => Kernel_inst_rematch000_taxi_out_cmd_ready,
      rematch000_taxi_out_cmd_firstIdx => Kernel_inst_rematch000_taxi_out_cmd_firstIdx,
      rematch000_taxi_out_cmd_lastIdx  => Kernel_inst_rematch000_taxi_out_cmd_lastIdx,
      rematch000_taxi_out_cmd_tag      => Kernel_inst_rematch000_taxi_out_cmd_tag,
      rematch001_taxi_out_valid        => Kernel_inst_rematch001_taxi_out_valid,
      rematch001_taxi_out_ready        => Kernel_inst_rematch001_taxi_out_ready,
      rematch001_taxi_out_dvalid       => Kernel_inst_rematch001_taxi_out_dvalid,
      rematch001_taxi_out_last         => Kernel_inst_rematch001_taxi_out_last,
      rematch001_taxi_out              => Kernel_inst_rematch001_taxi_out,
      rematch001_taxi_out_unl_valid    => Kernel_inst_rematch001_taxi_out_unl_valid,
      rematch001_taxi_out_unl_ready    => Kernel_inst_rematch001_taxi_out_unl_ready,
      rematch001_taxi_out_unl_tag      => Kernel_inst_rematch001_taxi_out_unl_tag,
      rematch001_taxi_out_cmd_valid    => Kernel_inst_rematch001_taxi_out_cmd_valid,
      rematch001_taxi_out_cmd_ready    => Kernel_inst_rematch001_taxi_out_cmd_ready,
      rematch001_taxi_out_cmd_firstIdx => Kernel_inst_rematch001_taxi_out_cmd_firstIdx,
      rematch001_taxi_out_cmd_lastIdx  => Kernel_inst_rematch001_taxi_out_cmd_lastIdx,
      rematch001_taxi_out_cmd_tag      => Kernel_inst_rematch001_taxi_out_cmd_tag,
      rematch002_taxi_out_valid        => Kernel_inst_rematch002_taxi_out_valid,
      rematch002_taxi_out_ready        => Kernel_inst_rematch002_taxi_out_ready,
      rematch002_taxi_out_dvalid       => Kernel_inst_rematch002_taxi_out_dvalid,
      rematch002_taxi_out_last         => Kernel_inst_rematch002_taxi_out_last,
      rematch002_taxi_out              => Kernel_inst_rematch002_taxi_out,
      rematch002_taxi_out_unl_valid    => Kernel_inst_rematch002_taxi_out_unl_valid,
      rematch002_taxi_out_unl_ready    => Kernel_inst_rematch002_taxi_out_unl_ready,
      rematch002_taxi_out_unl_tag      => Kernel_inst_rematch002_taxi_out_unl_tag,
      rematch002_taxi_out_cmd_valid    => Kernel_inst_rematch002_taxi_out_cmd_valid,
      rematch002_taxi_out_cmd_ready    => Kernel_inst_rematch002_taxi_out_cmd_ready,
      rematch002_taxi_out_cmd_firstIdx => Kernel_inst_rematch002_taxi_out_cmd_firstIdx,
      rematch002_taxi_out_cmd_lastIdx  => Kernel_inst_rematch002_taxi_out_cmd_lastIdx,
      rematch002_taxi_out_cmd_tag      => Kernel_inst_rematch002_taxi_out_cmd_tag,
      rematch003_taxi_out_valid        => Kernel_inst_rematch003_taxi_out_valid,
      rematch003_taxi_out_ready        => Kernel_inst_rematch003_taxi_out_ready,
      rematch003_taxi_out_dvalid       => Kernel_inst_rematch003_taxi_out_dvalid,
      rematch003_taxi_out_last         => Kernel_inst_rematch003_taxi_out_last,
      rematch003_taxi_out              => Kernel_inst_rematch003_taxi_out,
      rematch003_taxi_out_unl_valid    => Kernel_inst_rematch003_taxi_out_unl_valid,
      rematch003_taxi_out_unl_ready    => Kernel_inst_rematch003_taxi_out_unl_ready,
      rematch003_taxi_out_unl_tag      => Kernel_inst_rematch003_taxi_out_unl_tag,
      rematch003_taxi_out_cmd_valid    => Kernel_inst_rematch003_taxi_out_cmd_valid,
      rematch003_taxi_out_cmd_ready    => Kernel_inst_rematch003_taxi_out_cmd_ready,
      rematch003_taxi_out_cmd_firstIdx => Kernel_inst_rematch003_taxi_out_cmd_firstIdx,
      rematch003_taxi_out_cmd_lastIdx  => Kernel_inst_rematch003_taxi_out_cmd_lastIdx,
      rematch003_taxi_out_cmd_tag      => Kernel_inst_rematch003_taxi_out_cmd_tag,
      rematch004_taxi_out_valid        => Kernel_inst_rematch004_taxi_out_valid,
      rematch004_taxi_out_ready        => Kernel_inst_rematch004_taxi_out_ready,
      rematch004_taxi_out_dvalid       => Kernel_inst_rematch004_taxi_out_dvalid,
      rematch004_taxi_out_last         => Kernel_inst_rematch004_taxi_out_last,
      rematch004_taxi_out              => Kernel_inst_rematch004_taxi_out,
      rematch004_taxi_out_unl_valid    => Kernel_inst_rematch004_taxi_out_unl_valid,
      rematch004_taxi_out_unl_ready    => Kernel_inst_rematch004_taxi_out_unl_ready,
      rematch004_taxi_out_unl_tag      => Kernel_inst_rematch004_taxi_out_unl_tag,
      rematch004_taxi_out_cmd_valid    => Kernel_inst_rematch004_taxi_out_cmd_valid,
      rematch004_taxi_out_cmd_ready    => Kernel_inst_rematch004_taxi_out_cmd_ready,
      rematch004_taxi_out_cmd_firstIdx => Kernel_inst_rematch004_taxi_out_cmd_firstIdx,
      rematch004_taxi_out_cmd_lastIdx  => Kernel_inst_rematch004_taxi_out_cmd_lastIdx,
      rematch004_taxi_out_cmd_tag      => Kernel_inst_rematch004_taxi_out_cmd_tag,
      rematch005_taxi_out_valid        => Kernel_inst_rematch005_taxi_out_valid,
      rematch005_taxi_out_ready        => Kernel_inst_rematch005_taxi_out_ready,
      rematch005_taxi_out_dvalid       => Kernel_inst_rematch005_taxi_out_dvalid,
      rematch005_taxi_out_last         => Kernel_inst_rematch005_taxi_out_last,
      rematch005_taxi_out              => Kernel_inst_rematch005_taxi_out,
      rematch005_taxi_out_unl_valid    => Kernel_inst_rematch005_taxi_out_unl_valid,
      rematch005_taxi_out_unl_ready    => Kernel_inst_rematch005_taxi_out_unl_ready,
      rematch005_taxi_out_unl_tag      => Kernel_inst_rematch005_taxi_out_unl_tag,
      rematch005_taxi_out_cmd_valid    => Kernel_inst_rematch005_taxi_out_cmd_valid,
      rematch005_taxi_out_cmd_ready    => Kernel_inst_rematch005_taxi_out_cmd_ready,
      rematch005_taxi_out_cmd_firstIdx => Kernel_inst_rematch005_taxi_out_cmd_firstIdx,
      rematch005_taxi_out_cmd_lastIdx  => Kernel_inst_rematch005_taxi_out_cmd_lastIdx,
      rematch005_taxi_out_cmd_tag      => Kernel_inst_rematch005_taxi_out_cmd_tag,
      rematch006_taxi_out_valid        => Kernel_inst_rematch006_taxi_out_valid,
      rematch006_taxi_out_ready        => Kernel_inst_rematch006_taxi_out_ready,
      rematch006_taxi_out_dvalid       => Kernel_inst_rematch006_taxi_out_dvalid,
      rematch006_taxi_out_last         => Kernel_inst_rematch006_taxi_out_last,
      rematch006_taxi_out              => Kernel_inst_rematch006_taxi_out,
      rematch006_taxi_out_unl_valid    => Kernel_inst_rematch006_taxi_out_unl_valid,
      rematch006_taxi_out_unl_ready    => Kernel_inst_rematch006_taxi_out_unl_ready,
      rematch006_taxi_out_unl_tag      => Kernel_inst_rematch006_taxi_out_unl_tag,
      rematch006_taxi_out_cmd_valid    => Kernel_inst_rematch006_taxi_out_cmd_valid,
      rematch006_taxi_out_cmd_ready    => Kernel_inst_rematch006_taxi_out_cmd_ready,
      rematch006_taxi_out_cmd_firstIdx => Kernel_inst_rematch006_taxi_out_cmd_firstIdx,
      rematch006_taxi_out_cmd_lastIdx  => Kernel_inst_rematch006_taxi_out_cmd_lastIdx,
      rematch006_taxi_out_cmd_tag      => Kernel_inst_rematch006_taxi_out_cmd_tag,
      rematch007_taxi_out_valid        => Kernel_inst_rematch007_taxi_out_valid,
      rematch007_taxi_out_ready        => Kernel_inst_rematch007_taxi_out_ready,
      rematch007_taxi_out_dvalid       => Kernel_inst_rematch007_taxi_out_dvalid,
      rematch007_taxi_out_last         => Kernel_inst_rematch007_taxi_out_last,
      rematch007_taxi_out              => Kernel_inst_rematch007_taxi_out,
      rematch007_taxi_out_unl_valid    => Kernel_inst_rematch007_taxi_out_unl_valid,
      rematch007_taxi_out_unl_ready    => Kernel_inst_rematch007_taxi_out_unl_ready,
      rematch007_taxi_out_unl_tag      => Kernel_inst_rematch007_taxi_out_unl_tag,
      rematch007_taxi_out_cmd_valid    => Kernel_inst_rematch007_taxi_out_cmd_valid,
      rematch007_taxi_out_cmd_ready    => Kernel_inst_rematch007_taxi_out_cmd_ready,
      rematch007_taxi_out_cmd_firstIdx => Kernel_inst_rematch007_taxi_out_cmd_firstIdx,
      rematch007_taxi_out_cmd_lastIdx  => Kernel_inst_rematch007_taxi_out_cmd_lastIdx,
      rematch007_taxi_out_cmd_tag      => Kernel_inst_rematch007_taxi_out_cmd_tag,
      rematch008_taxi_out_valid        => Kernel_inst_rematch008_taxi_out_valid,
      rematch008_taxi_out_ready        => Kernel_inst_rematch008_taxi_out_ready,
      rematch008_taxi_out_dvalid       => Kernel_inst_rematch008_taxi_out_dvalid,
      rematch008_taxi_out_last         => Kernel_inst_rematch008_taxi_out_last,
      rematch008_taxi_out              => Kernel_inst_rematch008_taxi_out,
      rematch008_taxi_out_unl_valid    => Kernel_inst_rematch008_taxi_out_unl_valid,
      rematch008_taxi_out_unl_ready    => Kernel_inst_rematch008_taxi_out_unl_ready,
      rematch008_taxi_out_unl_tag      => Kernel_inst_rematch008_taxi_out_unl_tag,
      rematch008_taxi_out_cmd_valid    => Kernel_inst_rematch008_taxi_out_cmd_valid,
      rematch008_taxi_out_cmd_ready    => Kernel_inst_rematch008_taxi_out_cmd_ready,
      rematch008_taxi_out_cmd_firstIdx => Kernel_inst_rematch008_taxi_out_cmd_firstIdx,
      rematch008_taxi_out_cmd_lastIdx  => Kernel_inst_rematch008_taxi_out_cmd_lastIdx,
      rematch008_taxi_out_cmd_tag      => Kernel_inst_rematch008_taxi_out_cmd_tag,
      rematch009_taxi_out_valid        => Kernel_inst_rematch009_taxi_out_valid,
      rematch009_taxi_out_ready        => Kernel_inst_rematch009_taxi_out_ready,
      rematch009_taxi_out_dvalid       => Kernel_inst_rematch009_taxi_out_dvalid,
      rematch009_taxi_out_last         => Kernel_inst_rematch009_taxi_out_last,
      rematch009_taxi_out              => Kernel_inst_rematch009_taxi_out,
      rematch009_taxi_out_unl_valid    => Kernel_inst_rematch009_taxi_out_unl_valid,
      rematch009_taxi_out_unl_ready    => Kernel_inst_rematch009_taxi_out_unl_ready,
      rematch009_taxi_out_unl_tag      => Kernel_inst_rematch009_taxi_out_unl_tag,
      rematch009_taxi_out_cmd_valid    => Kernel_inst_rematch009_taxi_out_cmd_valid,
      rematch009_taxi_out_cmd_ready    => Kernel_inst_rematch009_taxi_out_cmd_ready,
      rematch009_taxi_out_cmd_firstIdx => Kernel_inst_rematch009_taxi_out_cmd_firstIdx,
      rematch009_taxi_out_cmd_lastIdx  => Kernel_inst_rematch009_taxi_out_cmd_lastIdx,
      rematch009_taxi_out_cmd_tag      => Kernel_inst_rematch009_taxi_out_cmd_tag,
      rematch010_taxi_out_valid        => Kernel_inst_rematch010_taxi_out_valid,
      rematch010_taxi_out_ready        => Kernel_inst_rematch010_taxi_out_ready,
      rematch010_taxi_out_dvalid       => Kernel_inst_rematch010_taxi_out_dvalid,
      rematch010_taxi_out_last         => Kernel_inst_rematch010_taxi_out_last,
      rematch010_taxi_out              => Kernel_inst_rematch010_taxi_out,
      rematch010_taxi_out_unl_valid    => Kernel_inst_rematch010_taxi_out_unl_valid,
      rematch010_taxi_out_unl_ready    => Kernel_inst_rematch010_taxi_out_unl_ready,
      rematch010_taxi_out_unl_tag      => Kernel_inst_rematch010_taxi_out_unl_tag,
      rematch010_taxi_out_cmd_valid    => Kernel_inst_rematch010_taxi_out_cmd_valid,
      rematch010_taxi_out_cmd_ready    => Kernel_inst_rematch010_taxi_out_cmd_ready,
      rematch010_taxi_out_cmd_firstIdx => Kernel_inst_rematch010_taxi_out_cmd_firstIdx,
      rematch010_taxi_out_cmd_lastIdx  => Kernel_inst_rematch010_taxi_out_cmd_lastIdx,
      rematch010_taxi_out_cmd_tag      => Kernel_inst_rematch010_taxi_out_cmd_tag,
      rematch011_taxi_out_valid        => Kernel_inst_rematch011_taxi_out_valid,
      rematch011_taxi_out_ready        => Kernel_inst_rematch011_taxi_out_ready,
      rematch011_taxi_out_dvalid       => Kernel_inst_rematch011_taxi_out_dvalid,
      rematch011_taxi_out_last         => Kernel_inst_rematch011_taxi_out_last,
      rematch011_taxi_out              => Kernel_inst_rematch011_taxi_out,
      rematch011_taxi_out_unl_valid    => Kernel_inst_rematch011_taxi_out_unl_valid,
      rematch011_taxi_out_unl_ready    => Kernel_inst_rematch011_taxi_out_unl_ready,
      rematch011_taxi_out_unl_tag      => Kernel_inst_rematch011_taxi_out_unl_tag,
      rematch011_taxi_out_cmd_valid    => Kernel_inst_rematch011_taxi_out_cmd_valid,
      rematch011_taxi_out_cmd_ready    => Kernel_inst_rematch011_taxi_out_cmd_ready,
      rematch011_taxi_out_cmd_firstIdx => Kernel_inst_rematch011_taxi_out_cmd_firstIdx,
      rematch011_taxi_out_cmd_lastIdx  => Kernel_inst_rematch011_taxi_out_cmd_lastIdx,
      rematch011_taxi_out_cmd_tag      => Kernel_inst_rematch011_taxi_out_cmd_tag,
      rematch012_taxi_out_valid        => Kernel_inst_rematch012_taxi_out_valid,
      rematch012_taxi_out_ready        => Kernel_inst_rematch012_taxi_out_ready,
      rematch012_taxi_out_dvalid       => Kernel_inst_rematch012_taxi_out_dvalid,
      rematch012_taxi_out_last         => Kernel_inst_rematch012_taxi_out_last,
      rematch012_taxi_out              => Kernel_inst_rematch012_taxi_out,
      rematch012_taxi_out_unl_valid    => Kernel_inst_rematch012_taxi_out_unl_valid,
      rematch012_taxi_out_unl_ready    => Kernel_inst_rematch012_taxi_out_unl_ready,
      rematch012_taxi_out_unl_tag      => Kernel_inst_rematch012_taxi_out_unl_tag,
      rematch012_taxi_out_cmd_valid    => Kernel_inst_rematch012_taxi_out_cmd_valid,
      rematch012_taxi_out_cmd_ready    => Kernel_inst_rematch012_taxi_out_cmd_ready,
      rematch012_taxi_out_cmd_firstIdx => Kernel_inst_rematch012_taxi_out_cmd_firstIdx,
      rematch012_taxi_out_cmd_lastIdx  => Kernel_inst_rematch012_taxi_out_cmd_lastIdx,
      rematch012_taxi_out_cmd_tag      => Kernel_inst_rematch012_taxi_out_cmd_tag,
      rematch013_taxi_out_valid        => Kernel_inst_rematch013_taxi_out_valid,
      rematch013_taxi_out_ready        => Kernel_inst_rematch013_taxi_out_ready,
      rematch013_taxi_out_dvalid       => Kernel_inst_rematch013_taxi_out_dvalid,
      rematch013_taxi_out_last         => Kernel_inst_rematch013_taxi_out_last,
      rematch013_taxi_out              => Kernel_inst_rematch013_taxi_out,
      rematch013_taxi_out_unl_valid    => Kernel_inst_rematch013_taxi_out_unl_valid,
      rematch013_taxi_out_unl_ready    => Kernel_inst_rematch013_taxi_out_unl_ready,
      rematch013_taxi_out_unl_tag      => Kernel_inst_rematch013_taxi_out_unl_tag,
      rematch013_taxi_out_cmd_valid    => Kernel_inst_rematch013_taxi_out_cmd_valid,
      rematch013_taxi_out_cmd_ready    => Kernel_inst_rematch013_taxi_out_cmd_ready,
      rematch013_taxi_out_cmd_firstIdx => Kernel_inst_rematch013_taxi_out_cmd_firstIdx,
      rematch013_taxi_out_cmd_lastIdx  => Kernel_inst_rematch013_taxi_out_cmd_lastIdx,
      rematch013_taxi_out_cmd_tag      => Kernel_inst_rematch013_taxi_out_cmd_tag,
      rematch014_taxi_out_valid        => Kernel_inst_rematch014_taxi_out_valid,
      rematch014_taxi_out_ready        => Kernel_inst_rematch014_taxi_out_ready,
      rematch014_taxi_out_dvalid       => Kernel_inst_rematch014_taxi_out_dvalid,
      rematch014_taxi_out_last         => Kernel_inst_rematch014_taxi_out_last,
      rematch014_taxi_out              => Kernel_inst_rematch014_taxi_out,
      rematch014_taxi_out_unl_valid    => Kernel_inst_rematch014_taxi_out_unl_valid,
      rematch014_taxi_out_unl_ready    => Kernel_inst_rematch014_taxi_out_unl_ready,
      rematch014_taxi_out_unl_tag      => Kernel_inst_rematch014_taxi_out_unl_tag,
      rematch014_taxi_out_cmd_valid    => Kernel_inst_rematch014_taxi_out_cmd_valid,
      rematch014_taxi_out_cmd_ready    => Kernel_inst_rematch014_taxi_out_cmd_ready,
      rematch014_taxi_out_cmd_firstIdx => Kernel_inst_rematch014_taxi_out_cmd_firstIdx,
      rematch014_taxi_out_cmd_lastIdx  => Kernel_inst_rematch014_taxi_out_cmd_lastIdx,
      rematch014_taxi_out_cmd_tag      => Kernel_inst_rematch014_taxi_out_cmd_tag,
      rematch015_taxi_out_valid        => Kernel_inst_rematch015_taxi_out_valid,
      rematch015_taxi_out_ready        => Kernel_inst_rematch015_taxi_out_ready,
      rematch015_taxi_out_dvalid       => Kernel_inst_rematch015_taxi_out_dvalid,
      rematch015_taxi_out_last         => Kernel_inst_rematch015_taxi_out_last,
      rematch015_taxi_out              => Kernel_inst_rematch015_taxi_out,
      rematch015_taxi_out_unl_valid    => Kernel_inst_rematch015_taxi_out_unl_valid,
      rematch015_taxi_out_unl_ready    => Kernel_inst_rematch015_taxi_out_unl_ready,
      rematch015_taxi_out_unl_tag      => Kernel_inst_rematch015_taxi_out_unl_tag,
      rematch015_taxi_out_cmd_valid    => Kernel_inst_rematch015_taxi_out_cmd_valid,
      rematch015_taxi_out_cmd_ready    => Kernel_inst_rematch015_taxi_out_cmd_ready,
      rematch015_taxi_out_cmd_firstIdx => Kernel_inst_rematch015_taxi_out_cmd_firstIdx,
      rematch015_taxi_out_cmd_lastIdx  => Kernel_inst_rematch015_taxi_out_cmd_lastIdx,
      rematch015_taxi_out_cmd_tag      => Kernel_inst_rematch015_taxi_out_cmd_tag,
      start                            => Kernel_inst_start,
      stop                             => Kernel_inst_stop,
      reset                            => Kernel_inst_reset,
      idle                             => Kernel_inst_idle,
      busy                             => Kernel_inst_busy,
      done                             => Kernel_inst_done,
      result                           => Kernel_inst_result,
      rematch000_firstidx              => Kernel_inst_rematch000_firstidx,
      rematch000_lastidx               => Kernel_inst_rematch000_lastidx,
      rematch001_firstidx              => Kernel_inst_rematch001_firstidx,
      rematch001_lastidx               => Kernel_inst_rematch001_lastidx,
      rematch002_firstidx              => Kernel_inst_rematch002_firstidx,
      rematch002_lastidx               => Kernel_inst_rematch002_lastidx,
      rematch003_firstidx              => Kernel_inst_rematch003_firstidx,
      rematch003_lastidx               => Kernel_inst_rematch003_lastidx,
      rematch004_firstidx              => Kernel_inst_rematch004_firstidx,
      rematch004_lastidx               => Kernel_inst_rematch004_lastidx,
      rematch005_firstidx              => Kernel_inst_rematch005_firstidx,
      rematch005_lastidx               => Kernel_inst_rematch005_lastidx,
      rematch006_firstidx              => Kernel_inst_rematch006_firstidx,
      rematch006_lastidx               => Kernel_inst_rematch006_lastidx,
      rematch007_firstidx              => Kernel_inst_rematch007_firstidx,
      rematch007_lastidx               => Kernel_inst_rematch007_lastidx,
      rematch008_firstidx              => Kernel_inst_rematch008_firstidx,
      rematch008_lastidx               => Kernel_inst_rematch008_lastidx,
      rematch009_firstidx              => Kernel_inst_rematch009_firstidx,
      rematch009_lastidx               => Kernel_inst_rematch009_lastidx,
      rematch010_firstidx              => Kernel_inst_rematch010_firstidx,
      rematch010_lastidx               => Kernel_inst_rematch010_lastidx,
      rematch011_firstidx              => Kernel_inst_rematch011_firstidx,
      rematch011_lastidx               => Kernel_inst_rematch011_lastidx,
      rematch012_firstidx              => Kernel_inst_rematch012_firstidx,
      rematch012_lastidx               => Kernel_inst_rematch012_lastidx,
      rematch013_firstidx              => Kernel_inst_rematch013_firstidx,
      rematch013_lastidx               => Kernel_inst_rematch013_lastidx,
      rematch014_firstidx              => Kernel_inst_rematch014_firstidx,
      rematch014_lastidx               => Kernel_inst_rematch014_lastidx,
      rematch015_firstidx              => Kernel_inst_rematch015_firstidx,
      rematch015_lastidx               => Kernel_inst_rematch015_lastidx,
      rematch000_taxi_firstidx         => Kernel_inst_rematch000_taxi_firstidx,
      rematch000_taxi_lastidx          => Kernel_inst_rematch000_taxi_lastidx,
      rematch001_taxi_firstidx         => Kernel_inst_rematch001_taxi_firstidx,
      rematch001_taxi_lastidx          => Kernel_inst_rematch001_taxi_lastidx,
      rematch002_taxi_firstidx         => Kernel_inst_rematch002_taxi_firstidx,
      rematch002_taxi_lastidx          => Kernel_inst_rematch002_taxi_lastidx,
      rematch003_taxi_firstidx         => Kernel_inst_rematch003_taxi_firstidx,
      rematch003_taxi_lastidx          => Kernel_inst_rematch003_taxi_lastidx,
      rematch004_taxi_firstidx         => Kernel_inst_rematch004_taxi_firstidx,
      rematch004_taxi_lastidx          => Kernel_inst_rematch004_taxi_lastidx,
      rematch005_taxi_firstidx         => Kernel_inst_rematch005_taxi_firstidx,
      rematch005_taxi_lastidx          => Kernel_inst_rematch005_taxi_lastidx,
      rematch006_taxi_firstidx         => Kernel_inst_rematch006_taxi_firstidx,
      rematch006_taxi_lastidx          => Kernel_inst_rematch006_taxi_lastidx,
      rematch007_taxi_firstidx         => Kernel_inst_rematch007_taxi_firstidx,
      rematch007_taxi_lastidx          => Kernel_inst_rematch007_taxi_lastidx,
      rematch008_taxi_firstidx         => Kernel_inst_rematch008_taxi_firstidx,
      rematch008_taxi_lastidx          => Kernel_inst_rematch008_taxi_lastidx,
      rematch009_taxi_firstidx         => Kernel_inst_rematch009_taxi_firstidx,
      rematch009_taxi_lastidx          => Kernel_inst_rematch009_taxi_lastidx,
      rematch010_taxi_firstidx         => Kernel_inst_rematch010_taxi_firstidx,
      rematch010_taxi_lastidx          => Kernel_inst_rematch010_taxi_lastidx,
      rematch011_taxi_firstidx         => Kernel_inst_rematch011_taxi_firstidx,
      rematch011_taxi_lastidx          => Kernel_inst_rematch011_taxi_lastidx,
      rematch012_taxi_firstidx         => Kernel_inst_rematch012_taxi_firstidx,
      rematch012_taxi_lastidx          => Kernel_inst_rematch012_taxi_lastidx,
      rematch013_taxi_firstidx         => Kernel_inst_rematch013_taxi_firstidx,
      rematch013_taxi_lastidx          => Kernel_inst_rematch013_taxi_lastidx,
      rematch014_taxi_firstidx         => Kernel_inst_rematch014_taxi_firstidx,
      rematch014_taxi_lastidx          => Kernel_inst_rematch014_taxi_lastidx,
      rematch015_taxi_firstidx         => Kernel_inst_rematch015_taxi_firstidx,
      rematch015_taxi_lastidx          => Kernel_inst_rematch015_taxi_lastidx,
      rematch000_taxi_count            => Kernel_inst_rematch000_taxi_count,
      rematch000_errors                => Kernel_inst_rematch000_errors,
      rematch001_taxi_count            => Kernel_inst_rematch001_taxi_count,
      rematch001_errors                => Kernel_inst_rematch001_errors,
      rematch002_taxi_count            => Kernel_inst_rematch002_taxi_count,
      rematch002_errors                => Kernel_inst_rematch002_errors,
      rematch003_taxi_count            => Kernel_inst_rematch003_taxi_count,
      rematch003_errors                => Kernel_inst_rematch003_errors,
      rematch004_taxi_count            => Kernel_inst_rematch004_taxi_count,
      rematch004_errors                => Kernel_inst_rematch004_errors,
      rematch005_taxi_count            => Kernel_inst_rematch005_taxi_count,
      rematch005_errors                => Kernel_inst_rematch005_errors,
      rematch006_taxi_count            => Kernel_inst_rematch006_taxi_count,
      rematch006_errors                => Kernel_inst_rematch006_errors,
      rematch007_taxi_count            => Kernel_inst_rematch007_taxi_count,
      rematch007_errors                => Kernel_inst_rematch007_errors,
      rematch008_taxi_count            => Kernel_inst_rematch008_taxi_count,
      rematch008_errors                => Kernel_inst_rematch008_errors,
      rematch009_taxi_count            => Kernel_inst_rematch009_taxi_count,
      rematch009_errors                => Kernel_inst_rematch009_errors,
      rematch010_taxi_count            => Kernel_inst_rematch010_taxi_count,
      rematch010_errors                => Kernel_inst_rematch010_errors,
      rematch011_taxi_count            => Kernel_inst_rematch011_taxi_count,
      rematch011_errors                => Kernel_inst_rematch011_errors,
      rematch012_taxi_count            => Kernel_inst_rematch012_taxi_count,
      rematch012_errors                => Kernel_inst_rematch012_errors,
      rematch013_taxi_count            => Kernel_inst_rematch013_taxi_count,
      rematch013_errors                => Kernel_inst_rematch013_errors,
      rematch014_taxi_count            => Kernel_inst_rematch014_taxi_count,
      rematch014_errors                => Kernel_inst_rematch014_errors,
      rematch015_taxi_count            => Kernel_inst_rematch015_taxi_count,
      rematch015_errors                => Kernel_inst_rematch015_errors
    );

  mmio_inst : mmio
    port map (
      kcd_clk                            => kcd_clk,
      kcd_reset                          => kcd_reset,
      f_start_data                       => mmio_inst_f_start_data,
      f_stop_data                        => mmio_inst_f_stop_data,
      f_reset_data                       => mmio_inst_f_reset_data,
      f_idle_write_data                  => mmio_inst_f_idle_write_data,
      f_busy_write_data                  => mmio_inst_f_busy_write_data,
      f_done_write_data                  => mmio_inst_f_done_write_data,
      f_result_write_data                => mmio_inst_f_result_write_data,
      f_rematch000_firstidx_data         => mmio_inst_f_rematch000_firstidx_data,
      f_rematch000_lastidx_data          => mmio_inst_f_rematch000_lastidx_data,
      f_rematch001_firstidx_data         => mmio_inst_f_rematch001_firstidx_data,
      f_rematch001_lastidx_data          => mmio_inst_f_rematch001_lastidx_data,
      f_rematch002_firstidx_data         => mmio_inst_f_rematch002_firstidx_data,
      f_rematch002_lastidx_data          => mmio_inst_f_rematch002_lastidx_data,
      f_rematch003_firstidx_data         => mmio_inst_f_rematch003_firstidx_data,
      f_rematch003_lastidx_data          => mmio_inst_f_rematch003_lastidx_data,
      f_rematch004_firstidx_data         => mmio_inst_f_rematch004_firstidx_data,
      f_rematch004_lastidx_data          => mmio_inst_f_rematch004_lastidx_data,
      f_rematch005_firstidx_data         => mmio_inst_f_rematch005_firstidx_data,
      f_rematch005_lastidx_data          => mmio_inst_f_rematch005_lastidx_data,
      f_rematch006_firstidx_data         => mmio_inst_f_rematch006_firstidx_data,
      f_rematch006_lastidx_data          => mmio_inst_f_rematch006_lastidx_data,
      f_rematch007_firstidx_data         => mmio_inst_f_rematch007_firstidx_data,
      f_rematch007_lastidx_data          => mmio_inst_f_rematch007_lastidx_data,
      f_rematch008_firstidx_data         => mmio_inst_f_rematch008_firstidx_data,
      f_rematch008_lastidx_data          => mmio_inst_f_rematch008_lastidx_data,
      f_rematch009_firstidx_data         => mmio_inst_f_rematch009_firstidx_data,
      f_rematch009_lastidx_data          => mmio_inst_f_rematch009_lastidx_data,
      f_rematch010_firstidx_data         => mmio_inst_f_rematch010_firstidx_data,
      f_rematch010_lastidx_data          => mmio_inst_f_rematch010_lastidx_data,
      f_rematch011_firstidx_data         => mmio_inst_f_rematch011_firstidx_data,
      f_rematch011_lastidx_data          => mmio_inst_f_rematch011_lastidx_data,
      f_rematch012_firstidx_data         => mmio_inst_f_rematch012_firstidx_data,
      f_rematch012_lastidx_data          => mmio_inst_f_rematch012_lastidx_data,
      f_rematch013_firstidx_data         => mmio_inst_f_rematch013_firstidx_data,
      f_rematch013_lastidx_data          => mmio_inst_f_rematch013_lastidx_data,
      f_rematch014_firstidx_data         => mmio_inst_f_rematch014_firstidx_data,
      f_rematch014_lastidx_data          => mmio_inst_f_rematch014_lastidx_data,
      f_rematch015_firstidx_data         => mmio_inst_f_rematch015_firstidx_data,
      f_rematch015_lastidx_data          => mmio_inst_f_rematch015_lastidx_data,
      f_rematch000_taxi_firstidx_data    => mmio_inst_f_rematch000_taxi_firstidx_data,
      f_rematch000_taxi_lastidx_data     => mmio_inst_f_rematch000_taxi_lastidx_data,
      f_rematch001_taxi_firstidx_data    => mmio_inst_f_rematch001_taxi_firstidx_data,
      f_rematch001_taxi_lastidx_data     => mmio_inst_f_rematch001_taxi_lastidx_data,
      f_rematch002_taxi_firstidx_data    => mmio_inst_f_rematch002_taxi_firstidx_data,
      f_rematch002_taxi_lastidx_data     => mmio_inst_f_rematch002_taxi_lastidx_data,
      f_rematch003_taxi_firstidx_data    => mmio_inst_f_rematch003_taxi_firstidx_data,
      f_rematch003_taxi_lastidx_data     => mmio_inst_f_rematch003_taxi_lastidx_data,
      f_rematch004_taxi_firstidx_data    => mmio_inst_f_rematch004_taxi_firstidx_data,
      f_rematch004_taxi_lastidx_data     => mmio_inst_f_rematch004_taxi_lastidx_data,
      f_rematch005_taxi_firstidx_data    => mmio_inst_f_rematch005_taxi_firstidx_data,
      f_rematch005_taxi_lastidx_data     => mmio_inst_f_rematch005_taxi_lastidx_data,
      f_rematch006_taxi_firstidx_data    => mmio_inst_f_rematch006_taxi_firstidx_data,
      f_rematch006_taxi_lastidx_data     => mmio_inst_f_rematch006_taxi_lastidx_data,
      f_rematch007_taxi_firstidx_data    => mmio_inst_f_rematch007_taxi_firstidx_data,
      f_rematch007_taxi_lastidx_data     => mmio_inst_f_rematch007_taxi_lastidx_data,
      f_rematch008_taxi_firstidx_data    => mmio_inst_f_rematch008_taxi_firstidx_data,
      f_rematch008_taxi_lastidx_data     => mmio_inst_f_rematch008_taxi_lastidx_data,
      f_rematch009_taxi_firstidx_data    => mmio_inst_f_rematch009_taxi_firstidx_data,
      f_rematch009_taxi_lastidx_data     => mmio_inst_f_rematch009_taxi_lastidx_data,
      f_rematch010_taxi_firstidx_data    => mmio_inst_f_rematch010_taxi_firstidx_data,
      f_rematch010_taxi_lastidx_data     => mmio_inst_f_rematch010_taxi_lastidx_data,
      f_rematch011_taxi_firstidx_data    => mmio_inst_f_rematch011_taxi_firstidx_data,
      f_rematch011_taxi_lastidx_data     => mmio_inst_f_rematch011_taxi_lastidx_data,
      f_rematch012_taxi_firstidx_data    => mmio_inst_f_rematch012_taxi_firstidx_data,
      f_rematch012_taxi_lastidx_data     => mmio_inst_f_rematch012_taxi_lastidx_data,
      f_rematch013_taxi_firstidx_data    => mmio_inst_f_rematch013_taxi_firstidx_data,
      f_rematch013_taxi_lastidx_data     => mmio_inst_f_rematch013_taxi_lastidx_data,
      f_rematch014_taxi_firstidx_data    => mmio_inst_f_rematch014_taxi_firstidx_data,
      f_rematch014_taxi_lastidx_data     => mmio_inst_f_rematch014_taxi_lastidx_data,
      f_rematch015_taxi_firstidx_data    => mmio_inst_f_rematch015_taxi_firstidx_data,
      f_rematch015_taxi_lastidx_data     => mmio_inst_f_rematch015_taxi_lastidx_data,
      f_rematch000_in_offsets_data       => mmio_inst_f_rematch000_in_offsets_data,
      f_rematch000_in_values_data        => mmio_inst_f_rematch000_in_values_data,
      f_rematch001_in_offsets_data       => mmio_inst_f_rematch001_in_offsets_data,
      f_rematch001_in_values_data        => mmio_inst_f_rematch001_in_values_data,
      f_rematch002_in_offsets_data       => mmio_inst_f_rematch002_in_offsets_data,
      f_rematch002_in_values_data        => mmio_inst_f_rematch002_in_values_data,
      f_rematch003_in_offsets_data       => mmio_inst_f_rematch003_in_offsets_data,
      f_rematch003_in_values_data        => mmio_inst_f_rematch003_in_values_data,
      f_rematch004_in_offsets_data       => mmio_inst_f_rematch004_in_offsets_data,
      f_rematch004_in_values_data        => mmio_inst_f_rematch004_in_values_data,
      f_rematch005_in_offsets_data       => mmio_inst_f_rematch005_in_offsets_data,
      f_rematch005_in_values_data        => mmio_inst_f_rematch005_in_values_data,
      f_rematch006_in_offsets_data       => mmio_inst_f_rematch006_in_offsets_data,
      f_rematch006_in_values_data        => mmio_inst_f_rematch006_in_values_data,
      f_rematch007_in_offsets_data       => mmio_inst_f_rematch007_in_offsets_data,
      f_rematch007_in_values_data        => mmio_inst_f_rematch007_in_values_data,
      f_rematch008_in_offsets_data       => mmio_inst_f_rematch008_in_offsets_data,
      f_rematch008_in_values_data        => mmio_inst_f_rematch008_in_values_data,
      f_rematch009_in_offsets_data       => mmio_inst_f_rematch009_in_offsets_data,
      f_rematch009_in_values_data        => mmio_inst_f_rematch009_in_values_data,
      f_rematch010_in_offsets_data       => mmio_inst_f_rematch010_in_offsets_data,
      f_rematch010_in_values_data        => mmio_inst_f_rematch010_in_values_data,
      f_rematch011_in_offsets_data       => mmio_inst_f_rematch011_in_offsets_data,
      f_rematch011_in_values_data        => mmio_inst_f_rematch011_in_values_data,
      f_rematch012_in_offsets_data       => mmio_inst_f_rematch012_in_offsets_data,
      f_rematch012_in_values_data        => mmio_inst_f_rematch012_in_values_data,
      f_rematch013_in_offsets_data       => mmio_inst_f_rematch013_in_offsets_data,
      f_rematch013_in_values_data        => mmio_inst_f_rematch013_in_values_data,
      f_rematch014_in_offsets_data       => mmio_inst_f_rematch014_in_offsets_data,
      f_rematch014_in_values_data        => mmio_inst_f_rematch014_in_values_data,
      f_rematch015_in_offsets_data       => mmio_inst_f_rematch015_in_offsets_data,
      f_rematch015_in_values_data        => mmio_inst_f_rematch015_in_values_data,
      f_rematch000_taxi_out_values_data  => mmio_inst_f_rematch000_taxi_out_values_data,
      f_rematch001_taxi_out_values_data  => mmio_inst_f_rematch001_taxi_out_values_data,
      f_rematch002_taxi_out_values_data  => mmio_inst_f_rematch002_taxi_out_values_data,
      f_rematch003_taxi_out_values_data  => mmio_inst_f_rematch003_taxi_out_values_data,
      f_rematch004_taxi_out_values_data  => mmio_inst_f_rematch004_taxi_out_values_data,
      f_rematch005_taxi_out_values_data  => mmio_inst_f_rematch005_taxi_out_values_data,
      f_rematch006_taxi_out_values_data  => mmio_inst_f_rematch006_taxi_out_values_data,
      f_rematch007_taxi_out_values_data  => mmio_inst_f_rematch007_taxi_out_values_data,
      f_rematch008_taxi_out_values_data  => mmio_inst_f_rematch008_taxi_out_values_data,
      f_rematch009_taxi_out_values_data  => mmio_inst_f_rematch009_taxi_out_values_data,
      f_rematch010_taxi_out_values_data  => mmio_inst_f_rematch010_taxi_out_values_data,
      f_rematch011_taxi_out_values_data  => mmio_inst_f_rematch011_taxi_out_values_data,
      f_rematch012_taxi_out_values_data  => mmio_inst_f_rematch012_taxi_out_values_data,
      f_rematch013_taxi_out_values_data  => mmio_inst_f_rematch013_taxi_out_values_data,
      f_rematch014_taxi_out_values_data  => mmio_inst_f_rematch014_taxi_out_values_data,
      f_rematch015_taxi_out_values_data  => mmio_inst_f_rematch015_taxi_out_values_data,
      f_rematch000_taxi_count_write_data => mmio_inst_f_rematch000_taxi_count_write_data,
      f_rematch000_errors_write_data     => mmio_inst_f_rematch000_errors_write_data,
      f_rematch001_taxi_count_write_data => mmio_inst_f_rematch001_taxi_count_write_data,
      f_rematch001_errors_write_data     => mmio_inst_f_rematch001_errors_write_data,
      f_rematch002_taxi_count_write_data => mmio_inst_f_rematch002_taxi_count_write_data,
      f_rematch002_errors_write_data     => mmio_inst_f_rematch002_errors_write_data,
      f_rematch003_taxi_count_write_data => mmio_inst_f_rematch003_taxi_count_write_data,
      f_rematch003_errors_write_data     => mmio_inst_f_rematch003_errors_write_data,
      f_rematch004_taxi_count_write_data => mmio_inst_f_rematch004_taxi_count_write_data,
      f_rematch004_errors_write_data     => mmio_inst_f_rematch004_errors_write_data,
      f_rematch005_taxi_count_write_data => mmio_inst_f_rematch005_taxi_count_write_data,
      f_rematch005_errors_write_data     => mmio_inst_f_rematch005_errors_write_data,
      f_rematch006_taxi_count_write_data => mmio_inst_f_rematch006_taxi_count_write_data,
      f_rematch006_errors_write_data     => mmio_inst_f_rematch006_errors_write_data,
      f_rematch007_taxi_count_write_data => mmio_inst_f_rematch007_taxi_count_write_data,
      f_rematch007_errors_write_data     => mmio_inst_f_rematch007_errors_write_data,
      f_rematch008_taxi_count_write_data => mmio_inst_f_rematch008_taxi_count_write_data,
      f_rematch008_errors_write_data     => mmio_inst_f_rematch008_errors_write_data,
      f_rematch009_taxi_count_write_data => mmio_inst_f_rematch009_taxi_count_write_data,
      f_rematch009_errors_write_data     => mmio_inst_f_rematch009_errors_write_data,
      f_rematch010_taxi_count_write_data => mmio_inst_f_rematch010_taxi_count_write_data,
      f_rematch010_errors_write_data     => mmio_inst_f_rematch010_errors_write_data,
      f_rematch011_taxi_count_write_data => mmio_inst_f_rematch011_taxi_count_write_data,
      f_rematch011_errors_write_data     => mmio_inst_f_rematch011_errors_write_data,
      f_rematch012_taxi_count_write_data => mmio_inst_f_rematch012_taxi_count_write_data,
      f_rematch012_errors_write_data     => mmio_inst_f_rematch012_errors_write_data,
      f_rematch013_taxi_count_write_data => mmio_inst_f_rematch013_taxi_count_write_data,
      f_rematch013_errors_write_data     => mmio_inst_f_rematch013_errors_write_data,
      f_rematch014_taxi_count_write_data => mmio_inst_f_rematch014_taxi_count_write_data,
      f_rematch014_errors_write_data     => mmio_inst_f_rematch014_errors_write_data,
      f_rematch015_taxi_count_write_data => mmio_inst_f_rematch015_taxi_count_write_data,
      f_rematch015_errors_write_data     => mmio_inst_f_rematch015_errors_write_data,
      mmio_awvalid                       => mmio_inst_mmio_awvalid,
      mmio_awready                       => mmio_inst_mmio_awready,
      mmio_awaddr                        => mmio_inst_mmio_awaddr,
      mmio_wvalid                        => mmio_inst_mmio_wvalid,
      mmio_wready                        => mmio_inst_mmio_wready,
      mmio_wdata                         => mmio_inst_mmio_wdata,
      mmio_wstrb                         => mmio_inst_mmio_wstrb,
      mmio_bvalid                        => mmio_inst_mmio_bvalid,
      mmio_bready                        => mmio_inst_mmio_bready,
      mmio_bresp                         => mmio_inst_mmio_bresp,
      mmio_arvalid                       => mmio_inst_mmio_arvalid,
      mmio_arready                       => mmio_inst_mmio_arready,
      mmio_araddr                        => mmio_inst_mmio_araddr,
      mmio_rvalid                        => mmio_inst_mmio_rvalid,
      mmio_rready                        => mmio_inst_mmio_rready,
      mmio_rdata                         => mmio_inst_mmio_rdata,
      mmio_rresp                         => mmio_inst_mmio_rresp
    );

  rematch000_in_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 2,
      BUS_ADDR_WIDTH => REMATCH000_IN_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch000_in_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch000_in_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch000_in_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch000_in_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch000_in_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch000_in_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch000_in_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch000_in_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch000_in_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch000_in_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch000_in_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch000_in_cmd_accm_inst_ctrl
    );

  rematch001_in_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 2,
      BUS_ADDR_WIDTH => REMATCH001_IN_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch001_in_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch001_in_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch001_in_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch001_in_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch001_in_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch001_in_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch001_in_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch001_in_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch001_in_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch001_in_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch001_in_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch001_in_cmd_accm_inst_ctrl
    );

  rematch002_in_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 2,
      BUS_ADDR_WIDTH => REMATCH002_IN_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch002_in_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch002_in_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch002_in_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch002_in_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch002_in_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch002_in_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch002_in_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch002_in_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch002_in_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch002_in_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch002_in_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch002_in_cmd_accm_inst_ctrl
    );

  rematch003_in_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 2,
      BUS_ADDR_WIDTH => REMATCH003_IN_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch003_in_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch003_in_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch003_in_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch003_in_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch003_in_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch003_in_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch003_in_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch003_in_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch003_in_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch003_in_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch003_in_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch003_in_cmd_accm_inst_ctrl
    );

  rematch004_in_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 2,
      BUS_ADDR_WIDTH => REMATCH004_IN_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch004_in_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch004_in_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch004_in_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch004_in_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch004_in_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch004_in_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch004_in_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch004_in_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch004_in_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch004_in_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch004_in_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch004_in_cmd_accm_inst_ctrl
    );

  rematch005_in_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 2,
      BUS_ADDR_WIDTH => REMATCH005_IN_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch005_in_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch005_in_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch005_in_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch005_in_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch005_in_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch005_in_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch005_in_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch005_in_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch005_in_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch005_in_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch005_in_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch005_in_cmd_accm_inst_ctrl
    );

  rematch006_in_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 2,
      BUS_ADDR_WIDTH => REMATCH006_IN_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch006_in_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch006_in_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch006_in_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch006_in_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch006_in_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch006_in_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch006_in_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch006_in_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch006_in_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch006_in_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch006_in_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch006_in_cmd_accm_inst_ctrl
    );

  rematch007_in_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 2,
      BUS_ADDR_WIDTH => REMATCH007_IN_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch007_in_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch007_in_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch007_in_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch007_in_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch007_in_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch007_in_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch007_in_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch007_in_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch007_in_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch007_in_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch007_in_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch007_in_cmd_accm_inst_ctrl
    );

  rematch008_in_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 2,
      BUS_ADDR_WIDTH => REMATCH008_IN_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch008_in_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch008_in_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch008_in_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch008_in_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch008_in_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch008_in_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch008_in_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch008_in_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch008_in_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch008_in_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch008_in_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch008_in_cmd_accm_inst_ctrl
    );

  rematch009_in_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 2,
      BUS_ADDR_WIDTH => REMATCH009_IN_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch009_in_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch009_in_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch009_in_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch009_in_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch009_in_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch009_in_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch009_in_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch009_in_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch009_in_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch009_in_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch009_in_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch009_in_cmd_accm_inst_ctrl
    );

  rematch010_in_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 2,
      BUS_ADDR_WIDTH => REMATCH010_IN_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch010_in_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch010_in_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch010_in_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch010_in_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch010_in_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch010_in_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch010_in_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch010_in_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch010_in_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch010_in_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch010_in_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch010_in_cmd_accm_inst_ctrl
    );

  rematch011_in_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 2,
      BUS_ADDR_WIDTH => REMATCH011_IN_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch011_in_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch011_in_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch011_in_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch011_in_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch011_in_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch011_in_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch011_in_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch011_in_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch011_in_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch011_in_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch011_in_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch011_in_cmd_accm_inst_ctrl
    );

  rematch012_in_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 2,
      BUS_ADDR_WIDTH => REMATCH012_IN_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch012_in_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch012_in_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch012_in_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch012_in_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch012_in_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch012_in_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch012_in_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch012_in_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch012_in_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch012_in_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch012_in_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch012_in_cmd_accm_inst_ctrl
    );

  rematch013_in_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 2,
      BUS_ADDR_WIDTH => REMATCH013_IN_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch013_in_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch013_in_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch013_in_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch013_in_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch013_in_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch013_in_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch013_in_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch013_in_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch013_in_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch013_in_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch013_in_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch013_in_cmd_accm_inst_ctrl
    );

  rematch014_in_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 2,
      BUS_ADDR_WIDTH => REMATCH014_IN_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch014_in_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch014_in_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch014_in_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch014_in_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch014_in_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch014_in_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch014_in_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch014_in_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch014_in_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch014_in_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch014_in_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch014_in_cmd_accm_inst_ctrl
    );

  rematch015_in_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 2,
      BUS_ADDR_WIDTH => REMATCH015_IN_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch015_in_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch015_in_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch015_in_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch015_in_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch015_in_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch015_in_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch015_in_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch015_in_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch015_in_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch015_in_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch015_in_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch015_in_cmd_accm_inst_ctrl
    );

  rematch000_taxi_out_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => REMATCH000_TAXI_OUT_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch000_taxi_out_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch000_taxi_out_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch000_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch000_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch000_taxi_out_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch000_taxi_out_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch000_taxi_out_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch000_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch000_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch000_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch000_taxi_out_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch000_taxi_out_cmd_accm_inst_ctrl
    );

  rematch001_taxi_out_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => REMATCH001_TAXI_OUT_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch001_taxi_out_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch001_taxi_out_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch001_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch001_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch001_taxi_out_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch001_taxi_out_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch001_taxi_out_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch001_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch001_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch001_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch001_taxi_out_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch001_taxi_out_cmd_accm_inst_ctrl
    );

  rematch002_taxi_out_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => REMATCH002_TAXI_OUT_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch002_taxi_out_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch002_taxi_out_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch002_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch002_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch002_taxi_out_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch002_taxi_out_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch002_taxi_out_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch002_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch002_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch002_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch002_taxi_out_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch002_taxi_out_cmd_accm_inst_ctrl
    );

  rematch003_taxi_out_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => REMATCH003_TAXI_OUT_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch003_taxi_out_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch003_taxi_out_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch003_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch003_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch003_taxi_out_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch003_taxi_out_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch003_taxi_out_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch003_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch003_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch003_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch003_taxi_out_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch003_taxi_out_cmd_accm_inst_ctrl
    );

  rematch004_taxi_out_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => REMATCH004_TAXI_OUT_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch004_taxi_out_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch004_taxi_out_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch004_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch004_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch004_taxi_out_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch004_taxi_out_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch004_taxi_out_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch004_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch004_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch004_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch004_taxi_out_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch004_taxi_out_cmd_accm_inst_ctrl
    );

  rematch005_taxi_out_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => REMATCH005_TAXI_OUT_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch005_taxi_out_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch005_taxi_out_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch005_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch005_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch005_taxi_out_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch005_taxi_out_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch005_taxi_out_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch005_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch005_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch005_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch005_taxi_out_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch005_taxi_out_cmd_accm_inst_ctrl
    );

  rematch006_taxi_out_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => REMATCH006_TAXI_OUT_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch006_taxi_out_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch006_taxi_out_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch006_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch006_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch006_taxi_out_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch006_taxi_out_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch006_taxi_out_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch006_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch006_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch006_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch006_taxi_out_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch006_taxi_out_cmd_accm_inst_ctrl
    );

  rematch007_taxi_out_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => REMATCH007_TAXI_OUT_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch007_taxi_out_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch007_taxi_out_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch007_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch007_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch007_taxi_out_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch007_taxi_out_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch007_taxi_out_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch007_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch007_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch007_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch007_taxi_out_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch007_taxi_out_cmd_accm_inst_ctrl
    );

  rematch008_taxi_out_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => REMATCH008_TAXI_OUT_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch008_taxi_out_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch008_taxi_out_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch008_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch008_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch008_taxi_out_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch008_taxi_out_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch008_taxi_out_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch008_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch008_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch008_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch008_taxi_out_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch008_taxi_out_cmd_accm_inst_ctrl
    );

  rematch009_taxi_out_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => REMATCH009_TAXI_OUT_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch009_taxi_out_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch009_taxi_out_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch009_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch009_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch009_taxi_out_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch009_taxi_out_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch009_taxi_out_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch009_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch009_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch009_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch009_taxi_out_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch009_taxi_out_cmd_accm_inst_ctrl
    );

  rematch010_taxi_out_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => REMATCH010_TAXI_OUT_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch010_taxi_out_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch010_taxi_out_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch010_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch010_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch010_taxi_out_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch010_taxi_out_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch010_taxi_out_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch010_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch010_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch010_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch010_taxi_out_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch010_taxi_out_cmd_accm_inst_ctrl
    );

  rematch011_taxi_out_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => REMATCH011_TAXI_OUT_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch011_taxi_out_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch011_taxi_out_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch011_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch011_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch011_taxi_out_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch011_taxi_out_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch011_taxi_out_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch011_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch011_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch011_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch011_taxi_out_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch011_taxi_out_cmd_accm_inst_ctrl
    );

  rematch012_taxi_out_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => REMATCH012_TAXI_OUT_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch012_taxi_out_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch012_taxi_out_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch012_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch012_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch012_taxi_out_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch012_taxi_out_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch012_taxi_out_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch012_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch012_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch012_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch012_taxi_out_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch012_taxi_out_cmd_accm_inst_ctrl
    );

  rematch013_taxi_out_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => REMATCH013_TAXI_OUT_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch013_taxi_out_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch013_taxi_out_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch013_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch013_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch013_taxi_out_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch013_taxi_out_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch013_taxi_out_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch013_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch013_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch013_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch013_taxi_out_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch013_taxi_out_cmd_accm_inst_ctrl
    );

  rematch014_taxi_out_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => REMATCH014_TAXI_OUT_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch014_taxi_out_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch014_taxi_out_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch014_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch014_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch014_taxi_out_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch014_taxi_out_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch014_taxi_out_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch014_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch014_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch014_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch014_taxi_out_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch014_taxi_out_cmd_accm_inst_ctrl
    );

  rematch015_taxi_out_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => REMATCH015_TAXI_OUT_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => rematch015_taxi_out_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => rematch015_taxi_out_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => rematch015_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => rematch015_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => rematch015_taxi_out_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => rematch015_taxi_out_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => rematch015_taxi_out_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => rematch015_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => rematch015_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => rematch015_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => rematch015_taxi_out_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => rematch015_taxi_out_cmd_accm_inst_ctrl
    );

  rematch000_in_cmd_valid                             <= rematch000_in_cmd_accm_inst_nucleus_cmd_valid;
  rematch000_in_cmd_accm_inst_nucleus_cmd_ready       <= rematch000_in_cmd_ready;
  rematch000_in_cmd_firstIdx                          <= rematch000_in_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch000_in_cmd_lastIdx                           <= rematch000_in_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch000_in_cmd_ctrl                              <= rematch000_in_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch000_in_cmd_tag                               <= rematch000_in_cmd_accm_inst_nucleus_cmd_tag;

  rematch001_in_cmd_valid                             <= rematch001_in_cmd_accm_inst_nucleus_cmd_valid;
  rematch001_in_cmd_accm_inst_nucleus_cmd_ready       <= rematch001_in_cmd_ready;
  rematch001_in_cmd_firstIdx                          <= rematch001_in_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch001_in_cmd_lastIdx                           <= rematch001_in_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch001_in_cmd_ctrl                              <= rematch001_in_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch001_in_cmd_tag                               <= rematch001_in_cmd_accm_inst_nucleus_cmd_tag;

  rematch002_in_cmd_valid                             <= rematch002_in_cmd_accm_inst_nucleus_cmd_valid;
  rematch002_in_cmd_accm_inst_nucleus_cmd_ready       <= rematch002_in_cmd_ready;
  rematch002_in_cmd_firstIdx                          <= rematch002_in_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch002_in_cmd_lastIdx                           <= rematch002_in_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch002_in_cmd_ctrl                              <= rematch002_in_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch002_in_cmd_tag                               <= rematch002_in_cmd_accm_inst_nucleus_cmd_tag;

  rematch003_in_cmd_valid                             <= rematch003_in_cmd_accm_inst_nucleus_cmd_valid;
  rematch003_in_cmd_accm_inst_nucleus_cmd_ready       <= rematch003_in_cmd_ready;
  rematch003_in_cmd_firstIdx                          <= rematch003_in_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch003_in_cmd_lastIdx                           <= rematch003_in_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch003_in_cmd_ctrl                              <= rematch003_in_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch003_in_cmd_tag                               <= rematch003_in_cmd_accm_inst_nucleus_cmd_tag;

  rematch004_in_cmd_valid                             <= rematch004_in_cmd_accm_inst_nucleus_cmd_valid;
  rematch004_in_cmd_accm_inst_nucleus_cmd_ready       <= rematch004_in_cmd_ready;
  rematch004_in_cmd_firstIdx                          <= rematch004_in_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch004_in_cmd_lastIdx                           <= rematch004_in_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch004_in_cmd_ctrl                              <= rematch004_in_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch004_in_cmd_tag                               <= rematch004_in_cmd_accm_inst_nucleus_cmd_tag;

  rematch005_in_cmd_valid                             <= rematch005_in_cmd_accm_inst_nucleus_cmd_valid;
  rematch005_in_cmd_accm_inst_nucleus_cmd_ready       <= rematch005_in_cmd_ready;
  rematch005_in_cmd_firstIdx                          <= rematch005_in_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch005_in_cmd_lastIdx                           <= rematch005_in_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch005_in_cmd_ctrl                              <= rematch005_in_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch005_in_cmd_tag                               <= rematch005_in_cmd_accm_inst_nucleus_cmd_tag;

  rematch006_in_cmd_valid                             <= rematch006_in_cmd_accm_inst_nucleus_cmd_valid;
  rematch006_in_cmd_accm_inst_nucleus_cmd_ready       <= rematch006_in_cmd_ready;
  rematch006_in_cmd_firstIdx                          <= rematch006_in_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch006_in_cmd_lastIdx                           <= rematch006_in_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch006_in_cmd_ctrl                              <= rematch006_in_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch006_in_cmd_tag                               <= rematch006_in_cmd_accm_inst_nucleus_cmd_tag;

  rematch007_in_cmd_valid                             <= rematch007_in_cmd_accm_inst_nucleus_cmd_valid;
  rematch007_in_cmd_accm_inst_nucleus_cmd_ready       <= rematch007_in_cmd_ready;
  rematch007_in_cmd_firstIdx                          <= rematch007_in_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch007_in_cmd_lastIdx                           <= rematch007_in_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch007_in_cmd_ctrl                              <= rematch007_in_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch007_in_cmd_tag                               <= rematch007_in_cmd_accm_inst_nucleus_cmd_tag;

  rematch008_in_cmd_valid                             <= rematch008_in_cmd_accm_inst_nucleus_cmd_valid;
  rematch008_in_cmd_accm_inst_nucleus_cmd_ready       <= rematch008_in_cmd_ready;
  rematch008_in_cmd_firstIdx                          <= rematch008_in_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch008_in_cmd_lastIdx                           <= rematch008_in_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch008_in_cmd_ctrl                              <= rematch008_in_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch008_in_cmd_tag                               <= rematch008_in_cmd_accm_inst_nucleus_cmd_tag;

  rematch009_in_cmd_valid                             <= rematch009_in_cmd_accm_inst_nucleus_cmd_valid;
  rematch009_in_cmd_accm_inst_nucleus_cmd_ready       <= rematch009_in_cmd_ready;
  rematch009_in_cmd_firstIdx                          <= rematch009_in_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch009_in_cmd_lastIdx                           <= rematch009_in_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch009_in_cmd_ctrl                              <= rematch009_in_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch009_in_cmd_tag                               <= rematch009_in_cmd_accm_inst_nucleus_cmd_tag;

  rematch010_in_cmd_valid                             <= rematch010_in_cmd_accm_inst_nucleus_cmd_valid;
  rematch010_in_cmd_accm_inst_nucleus_cmd_ready       <= rematch010_in_cmd_ready;
  rematch010_in_cmd_firstIdx                          <= rematch010_in_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch010_in_cmd_lastIdx                           <= rematch010_in_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch010_in_cmd_ctrl                              <= rematch010_in_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch010_in_cmd_tag                               <= rematch010_in_cmd_accm_inst_nucleus_cmd_tag;

  rematch011_in_cmd_valid                             <= rematch011_in_cmd_accm_inst_nucleus_cmd_valid;
  rematch011_in_cmd_accm_inst_nucleus_cmd_ready       <= rematch011_in_cmd_ready;
  rematch011_in_cmd_firstIdx                          <= rematch011_in_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch011_in_cmd_lastIdx                           <= rematch011_in_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch011_in_cmd_ctrl                              <= rematch011_in_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch011_in_cmd_tag                               <= rematch011_in_cmd_accm_inst_nucleus_cmd_tag;

  rematch012_in_cmd_valid                             <= rematch012_in_cmd_accm_inst_nucleus_cmd_valid;
  rematch012_in_cmd_accm_inst_nucleus_cmd_ready       <= rematch012_in_cmd_ready;
  rematch012_in_cmd_firstIdx                          <= rematch012_in_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch012_in_cmd_lastIdx                           <= rematch012_in_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch012_in_cmd_ctrl                              <= rematch012_in_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch012_in_cmd_tag                               <= rematch012_in_cmd_accm_inst_nucleus_cmd_tag;

  rematch013_in_cmd_valid                             <= rematch013_in_cmd_accm_inst_nucleus_cmd_valid;
  rematch013_in_cmd_accm_inst_nucleus_cmd_ready       <= rematch013_in_cmd_ready;
  rematch013_in_cmd_firstIdx                          <= rematch013_in_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch013_in_cmd_lastIdx                           <= rematch013_in_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch013_in_cmd_ctrl                              <= rematch013_in_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch013_in_cmd_tag                               <= rematch013_in_cmd_accm_inst_nucleus_cmd_tag;

  rematch014_in_cmd_valid                             <= rematch014_in_cmd_accm_inst_nucleus_cmd_valid;
  rematch014_in_cmd_accm_inst_nucleus_cmd_ready       <= rematch014_in_cmd_ready;
  rematch014_in_cmd_firstIdx                          <= rematch014_in_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch014_in_cmd_lastIdx                           <= rematch014_in_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch014_in_cmd_ctrl                              <= rematch014_in_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch014_in_cmd_tag                               <= rematch014_in_cmd_accm_inst_nucleus_cmd_tag;

  rematch015_in_cmd_valid                             <= rematch015_in_cmd_accm_inst_nucleus_cmd_valid;
  rematch015_in_cmd_accm_inst_nucleus_cmd_ready       <= rematch015_in_cmd_ready;
  rematch015_in_cmd_firstIdx                          <= rematch015_in_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch015_in_cmd_lastIdx                           <= rematch015_in_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch015_in_cmd_ctrl                              <= rematch015_in_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch015_in_cmd_tag                               <= rematch015_in_cmd_accm_inst_nucleus_cmd_tag;

  rematch000_taxi_out_valid                           <= Kernel_inst_rematch000_taxi_out_valid;
  Kernel_inst_rematch000_taxi_out_ready               <= rematch000_taxi_out_ready;
  rematch000_taxi_out_dvalid                          <= Kernel_inst_rematch000_taxi_out_dvalid;
  rematch000_taxi_out_last                            <= Kernel_inst_rematch000_taxi_out_last;
  rematch000_taxi_out                                 <= Kernel_inst_rematch000_taxi_out;

  rematch000_taxi_out_cmd_valid                       <= rematch000_taxi_out_cmd_accm_inst_nucleus_cmd_valid;
  rematch000_taxi_out_cmd_accm_inst_nucleus_cmd_ready <= rematch000_taxi_out_cmd_ready;
  rematch000_taxi_out_cmd_firstIdx                    <= rematch000_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch000_taxi_out_cmd_lastIdx                     <= rematch000_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch000_taxi_out_cmd_ctrl                        <= rematch000_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch000_taxi_out_cmd_tag                         <= rematch000_taxi_out_cmd_accm_inst_nucleus_cmd_tag;

  rematch001_taxi_out_valid                           <= Kernel_inst_rematch001_taxi_out_valid;
  Kernel_inst_rematch001_taxi_out_ready               <= rematch001_taxi_out_ready;
  rematch001_taxi_out_dvalid                          <= Kernel_inst_rematch001_taxi_out_dvalid;
  rematch001_taxi_out_last                            <= Kernel_inst_rematch001_taxi_out_last;
  rematch001_taxi_out                                 <= Kernel_inst_rematch001_taxi_out;

  rematch001_taxi_out_cmd_valid                       <= rematch001_taxi_out_cmd_accm_inst_nucleus_cmd_valid;
  rematch001_taxi_out_cmd_accm_inst_nucleus_cmd_ready <= rematch001_taxi_out_cmd_ready;
  rematch001_taxi_out_cmd_firstIdx                    <= rematch001_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch001_taxi_out_cmd_lastIdx                     <= rematch001_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch001_taxi_out_cmd_ctrl                        <= rematch001_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch001_taxi_out_cmd_tag                         <= rematch001_taxi_out_cmd_accm_inst_nucleus_cmd_tag;

  rematch002_taxi_out_valid                           <= Kernel_inst_rematch002_taxi_out_valid;
  Kernel_inst_rematch002_taxi_out_ready               <= rematch002_taxi_out_ready;
  rematch002_taxi_out_dvalid                          <= Kernel_inst_rematch002_taxi_out_dvalid;
  rematch002_taxi_out_last                            <= Kernel_inst_rematch002_taxi_out_last;
  rematch002_taxi_out                                 <= Kernel_inst_rematch002_taxi_out;

  rematch002_taxi_out_cmd_valid                       <= rematch002_taxi_out_cmd_accm_inst_nucleus_cmd_valid;
  rematch002_taxi_out_cmd_accm_inst_nucleus_cmd_ready <= rematch002_taxi_out_cmd_ready;
  rematch002_taxi_out_cmd_firstIdx                    <= rematch002_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch002_taxi_out_cmd_lastIdx                     <= rematch002_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch002_taxi_out_cmd_ctrl                        <= rematch002_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch002_taxi_out_cmd_tag                         <= rematch002_taxi_out_cmd_accm_inst_nucleus_cmd_tag;

  rematch003_taxi_out_valid                           <= Kernel_inst_rematch003_taxi_out_valid;
  Kernel_inst_rematch003_taxi_out_ready               <= rematch003_taxi_out_ready;
  rematch003_taxi_out_dvalid                          <= Kernel_inst_rematch003_taxi_out_dvalid;
  rematch003_taxi_out_last                            <= Kernel_inst_rematch003_taxi_out_last;
  rematch003_taxi_out                                 <= Kernel_inst_rematch003_taxi_out;

  rematch003_taxi_out_cmd_valid                       <= rematch003_taxi_out_cmd_accm_inst_nucleus_cmd_valid;
  rematch003_taxi_out_cmd_accm_inst_nucleus_cmd_ready <= rematch003_taxi_out_cmd_ready;
  rematch003_taxi_out_cmd_firstIdx                    <= rematch003_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch003_taxi_out_cmd_lastIdx                     <= rematch003_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch003_taxi_out_cmd_ctrl                        <= rematch003_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch003_taxi_out_cmd_tag                         <= rematch003_taxi_out_cmd_accm_inst_nucleus_cmd_tag;

  rematch004_taxi_out_valid                           <= Kernel_inst_rematch004_taxi_out_valid;
  Kernel_inst_rematch004_taxi_out_ready               <= rematch004_taxi_out_ready;
  rematch004_taxi_out_dvalid                          <= Kernel_inst_rematch004_taxi_out_dvalid;
  rematch004_taxi_out_last                            <= Kernel_inst_rematch004_taxi_out_last;
  rematch004_taxi_out                                 <= Kernel_inst_rematch004_taxi_out;

  rematch004_taxi_out_cmd_valid                       <= rematch004_taxi_out_cmd_accm_inst_nucleus_cmd_valid;
  rematch004_taxi_out_cmd_accm_inst_nucleus_cmd_ready <= rematch004_taxi_out_cmd_ready;
  rematch004_taxi_out_cmd_firstIdx                    <= rematch004_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch004_taxi_out_cmd_lastIdx                     <= rematch004_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch004_taxi_out_cmd_ctrl                        <= rematch004_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch004_taxi_out_cmd_tag                         <= rematch004_taxi_out_cmd_accm_inst_nucleus_cmd_tag;

  rematch005_taxi_out_valid                           <= Kernel_inst_rematch005_taxi_out_valid;
  Kernel_inst_rematch005_taxi_out_ready               <= rematch005_taxi_out_ready;
  rematch005_taxi_out_dvalid                          <= Kernel_inst_rematch005_taxi_out_dvalid;
  rematch005_taxi_out_last                            <= Kernel_inst_rematch005_taxi_out_last;
  rematch005_taxi_out                                 <= Kernel_inst_rematch005_taxi_out;

  rematch005_taxi_out_cmd_valid                       <= rematch005_taxi_out_cmd_accm_inst_nucleus_cmd_valid;
  rematch005_taxi_out_cmd_accm_inst_nucleus_cmd_ready <= rematch005_taxi_out_cmd_ready;
  rematch005_taxi_out_cmd_firstIdx                    <= rematch005_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch005_taxi_out_cmd_lastIdx                     <= rematch005_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch005_taxi_out_cmd_ctrl                        <= rematch005_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch005_taxi_out_cmd_tag                         <= rematch005_taxi_out_cmd_accm_inst_nucleus_cmd_tag;

  rematch006_taxi_out_valid                           <= Kernel_inst_rematch006_taxi_out_valid;
  Kernel_inst_rematch006_taxi_out_ready               <= rematch006_taxi_out_ready;
  rematch006_taxi_out_dvalid                          <= Kernel_inst_rematch006_taxi_out_dvalid;
  rematch006_taxi_out_last                            <= Kernel_inst_rematch006_taxi_out_last;
  rematch006_taxi_out                                 <= Kernel_inst_rematch006_taxi_out;

  rematch006_taxi_out_cmd_valid                       <= rematch006_taxi_out_cmd_accm_inst_nucleus_cmd_valid;
  rematch006_taxi_out_cmd_accm_inst_nucleus_cmd_ready <= rematch006_taxi_out_cmd_ready;
  rematch006_taxi_out_cmd_firstIdx                    <= rematch006_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch006_taxi_out_cmd_lastIdx                     <= rematch006_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch006_taxi_out_cmd_ctrl                        <= rematch006_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch006_taxi_out_cmd_tag                         <= rematch006_taxi_out_cmd_accm_inst_nucleus_cmd_tag;

  rematch007_taxi_out_valid                           <= Kernel_inst_rematch007_taxi_out_valid;
  Kernel_inst_rematch007_taxi_out_ready               <= rematch007_taxi_out_ready;
  rematch007_taxi_out_dvalid                          <= Kernel_inst_rematch007_taxi_out_dvalid;
  rematch007_taxi_out_last                            <= Kernel_inst_rematch007_taxi_out_last;
  rematch007_taxi_out                                 <= Kernel_inst_rematch007_taxi_out;

  rematch007_taxi_out_cmd_valid                       <= rematch007_taxi_out_cmd_accm_inst_nucleus_cmd_valid;
  rematch007_taxi_out_cmd_accm_inst_nucleus_cmd_ready <= rematch007_taxi_out_cmd_ready;
  rematch007_taxi_out_cmd_firstIdx                    <= rematch007_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch007_taxi_out_cmd_lastIdx                     <= rematch007_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch007_taxi_out_cmd_ctrl                        <= rematch007_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch007_taxi_out_cmd_tag                         <= rematch007_taxi_out_cmd_accm_inst_nucleus_cmd_tag;

  rematch008_taxi_out_valid                           <= Kernel_inst_rematch008_taxi_out_valid;
  Kernel_inst_rematch008_taxi_out_ready               <= rematch008_taxi_out_ready;
  rematch008_taxi_out_dvalid                          <= Kernel_inst_rematch008_taxi_out_dvalid;
  rematch008_taxi_out_last                            <= Kernel_inst_rematch008_taxi_out_last;
  rematch008_taxi_out                                 <= Kernel_inst_rematch008_taxi_out;

  rematch008_taxi_out_cmd_valid                       <= rematch008_taxi_out_cmd_accm_inst_nucleus_cmd_valid;
  rematch008_taxi_out_cmd_accm_inst_nucleus_cmd_ready <= rematch008_taxi_out_cmd_ready;
  rematch008_taxi_out_cmd_firstIdx                    <= rematch008_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch008_taxi_out_cmd_lastIdx                     <= rematch008_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch008_taxi_out_cmd_ctrl                        <= rematch008_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch008_taxi_out_cmd_tag                         <= rematch008_taxi_out_cmd_accm_inst_nucleus_cmd_tag;

  rematch009_taxi_out_valid                           <= Kernel_inst_rematch009_taxi_out_valid;
  Kernel_inst_rematch009_taxi_out_ready               <= rematch009_taxi_out_ready;
  rematch009_taxi_out_dvalid                          <= Kernel_inst_rematch009_taxi_out_dvalid;
  rematch009_taxi_out_last                            <= Kernel_inst_rematch009_taxi_out_last;
  rematch009_taxi_out                                 <= Kernel_inst_rematch009_taxi_out;

  rematch009_taxi_out_cmd_valid                       <= rematch009_taxi_out_cmd_accm_inst_nucleus_cmd_valid;
  rematch009_taxi_out_cmd_accm_inst_nucleus_cmd_ready <= rematch009_taxi_out_cmd_ready;
  rematch009_taxi_out_cmd_firstIdx                    <= rematch009_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch009_taxi_out_cmd_lastIdx                     <= rematch009_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch009_taxi_out_cmd_ctrl                        <= rematch009_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch009_taxi_out_cmd_tag                         <= rematch009_taxi_out_cmd_accm_inst_nucleus_cmd_tag;

  rematch010_taxi_out_valid                           <= Kernel_inst_rematch010_taxi_out_valid;
  Kernel_inst_rematch010_taxi_out_ready               <= rematch010_taxi_out_ready;
  rematch010_taxi_out_dvalid                          <= Kernel_inst_rematch010_taxi_out_dvalid;
  rematch010_taxi_out_last                            <= Kernel_inst_rematch010_taxi_out_last;
  rematch010_taxi_out                                 <= Kernel_inst_rematch010_taxi_out;

  rematch010_taxi_out_cmd_valid                       <= rematch010_taxi_out_cmd_accm_inst_nucleus_cmd_valid;
  rematch010_taxi_out_cmd_accm_inst_nucleus_cmd_ready <= rematch010_taxi_out_cmd_ready;
  rematch010_taxi_out_cmd_firstIdx                    <= rematch010_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch010_taxi_out_cmd_lastIdx                     <= rematch010_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch010_taxi_out_cmd_ctrl                        <= rematch010_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch010_taxi_out_cmd_tag                         <= rematch010_taxi_out_cmd_accm_inst_nucleus_cmd_tag;

  rematch011_taxi_out_valid                           <= Kernel_inst_rematch011_taxi_out_valid;
  Kernel_inst_rematch011_taxi_out_ready               <= rematch011_taxi_out_ready;
  rematch011_taxi_out_dvalid                          <= Kernel_inst_rematch011_taxi_out_dvalid;
  rematch011_taxi_out_last                            <= Kernel_inst_rematch011_taxi_out_last;
  rematch011_taxi_out                                 <= Kernel_inst_rematch011_taxi_out;

  rematch011_taxi_out_cmd_valid                       <= rematch011_taxi_out_cmd_accm_inst_nucleus_cmd_valid;
  rematch011_taxi_out_cmd_accm_inst_nucleus_cmd_ready <= rematch011_taxi_out_cmd_ready;
  rematch011_taxi_out_cmd_firstIdx                    <= rematch011_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch011_taxi_out_cmd_lastIdx                     <= rematch011_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch011_taxi_out_cmd_ctrl                        <= rematch011_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch011_taxi_out_cmd_tag                         <= rematch011_taxi_out_cmd_accm_inst_nucleus_cmd_tag;

  rematch012_taxi_out_valid                           <= Kernel_inst_rematch012_taxi_out_valid;
  Kernel_inst_rematch012_taxi_out_ready               <= rematch012_taxi_out_ready;
  rematch012_taxi_out_dvalid                          <= Kernel_inst_rematch012_taxi_out_dvalid;
  rematch012_taxi_out_last                            <= Kernel_inst_rematch012_taxi_out_last;
  rematch012_taxi_out                                 <= Kernel_inst_rematch012_taxi_out;

  rematch012_taxi_out_cmd_valid                       <= rematch012_taxi_out_cmd_accm_inst_nucleus_cmd_valid;
  rematch012_taxi_out_cmd_accm_inst_nucleus_cmd_ready <= rematch012_taxi_out_cmd_ready;
  rematch012_taxi_out_cmd_firstIdx                    <= rematch012_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch012_taxi_out_cmd_lastIdx                     <= rematch012_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch012_taxi_out_cmd_ctrl                        <= rematch012_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch012_taxi_out_cmd_tag                         <= rematch012_taxi_out_cmd_accm_inst_nucleus_cmd_tag;

  rematch013_taxi_out_valid                           <= Kernel_inst_rematch013_taxi_out_valid;
  Kernel_inst_rematch013_taxi_out_ready               <= rematch013_taxi_out_ready;
  rematch013_taxi_out_dvalid                          <= Kernel_inst_rematch013_taxi_out_dvalid;
  rematch013_taxi_out_last                            <= Kernel_inst_rematch013_taxi_out_last;
  rematch013_taxi_out                                 <= Kernel_inst_rematch013_taxi_out;

  rematch013_taxi_out_cmd_valid                       <= rematch013_taxi_out_cmd_accm_inst_nucleus_cmd_valid;
  rematch013_taxi_out_cmd_accm_inst_nucleus_cmd_ready <= rematch013_taxi_out_cmd_ready;
  rematch013_taxi_out_cmd_firstIdx                    <= rematch013_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch013_taxi_out_cmd_lastIdx                     <= rematch013_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch013_taxi_out_cmd_ctrl                        <= rematch013_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch013_taxi_out_cmd_tag                         <= rematch013_taxi_out_cmd_accm_inst_nucleus_cmd_tag;

  rematch014_taxi_out_valid                           <= Kernel_inst_rematch014_taxi_out_valid;
  Kernel_inst_rematch014_taxi_out_ready               <= rematch014_taxi_out_ready;
  rematch014_taxi_out_dvalid                          <= Kernel_inst_rematch014_taxi_out_dvalid;
  rematch014_taxi_out_last                            <= Kernel_inst_rematch014_taxi_out_last;
  rematch014_taxi_out                                 <= Kernel_inst_rematch014_taxi_out;

  rematch014_taxi_out_cmd_valid                       <= rematch014_taxi_out_cmd_accm_inst_nucleus_cmd_valid;
  rematch014_taxi_out_cmd_accm_inst_nucleus_cmd_ready <= rematch014_taxi_out_cmd_ready;
  rematch014_taxi_out_cmd_firstIdx                    <= rematch014_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch014_taxi_out_cmd_lastIdx                     <= rematch014_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch014_taxi_out_cmd_ctrl                        <= rematch014_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch014_taxi_out_cmd_tag                         <= rematch014_taxi_out_cmd_accm_inst_nucleus_cmd_tag;

  rematch015_taxi_out_valid                           <= Kernel_inst_rematch015_taxi_out_valid;
  Kernel_inst_rematch015_taxi_out_ready               <= rematch015_taxi_out_ready;
  rematch015_taxi_out_dvalid                          <= Kernel_inst_rematch015_taxi_out_dvalid;
  rematch015_taxi_out_last                            <= Kernel_inst_rematch015_taxi_out_last;
  rematch015_taxi_out                                 <= Kernel_inst_rematch015_taxi_out;

  rematch015_taxi_out_cmd_valid                       <= rematch015_taxi_out_cmd_accm_inst_nucleus_cmd_valid;
  rematch015_taxi_out_cmd_accm_inst_nucleus_cmd_ready <= rematch015_taxi_out_cmd_ready;
  rematch015_taxi_out_cmd_firstIdx                    <= rematch015_taxi_out_cmd_accm_inst_nucleus_cmd_firstIdx;
  rematch015_taxi_out_cmd_lastIdx                     <= rematch015_taxi_out_cmd_accm_inst_nucleus_cmd_lastIdx;
  rematch015_taxi_out_cmd_ctrl                        <= rematch015_taxi_out_cmd_accm_inst_nucleus_cmd_ctrl;
  rematch015_taxi_out_cmd_tag                         <= rematch015_taxi_out_cmd_accm_inst_nucleus_cmd_tag;

  Kernel_inst_rematch000_in_valid                       <= rematch000_in_valid;
  rematch000_in_ready                                   <= Kernel_inst_rematch000_in_ready;
  Kernel_inst_rematch000_in_dvalid                      <= rematch000_in_dvalid;
  Kernel_inst_rematch000_in_last                        <= rematch000_in_last;
  Kernel_inst_rematch000_in_length                      <= rematch000_in_length;
  Kernel_inst_rematch000_in_count                       <= rematch000_in_count;
  Kernel_inst_rematch000_in_chars_valid                 <= rematch000_in_chars_valid;
  rematch000_in_chars_ready                             <= Kernel_inst_rematch000_in_chars_ready;
  Kernel_inst_rematch000_in_chars_dvalid                <= rematch000_in_chars_dvalid;
  Kernel_inst_rematch000_in_chars_last                  <= rematch000_in_chars_last;
  Kernel_inst_rematch000_in_chars                       <= rematch000_in_chars;
  Kernel_inst_rematch000_in_chars_count                 <= rematch000_in_chars_count;

  Kernel_inst_rematch000_in_unl_valid                   <= rematch000_in_unl_valid;
  rematch000_in_unl_ready                               <= Kernel_inst_rematch000_in_unl_ready;
  Kernel_inst_rematch000_in_unl_tag                     <= rematch000_in_unl_tag;

  Kernel_inst_rematch001_in_valid                       <= rematch001_in_valid;
  rematch001_in_ready                                   <= Kernel_inst_rematch001_in_ready;
  Kernel_inst_rematch001_in_dvalid                      <= rematch001_in_dvalid;
  Kernel_inst_rematch001_in_last                        <= rematch001_in_last;
  Kernel_inst_rematch001_in_length                      <= rematch001_in_length;
  Kernel_inst_rematch001_in_count                       <= rematch001_in_count;
  Kernel_inst_rematch001_in_chars_valid                 <= rematch001_in_chars_valid;
  rematch001_in_chars_ready                             <= Kernel_inst_rematch001_in_chars_ready;
  Kernel_inst_rematch001_in_chars_dvalid                <= rematch001_in_chars_dvalid;
  Kernel_inst_rematch001_in_chars_last                  <= rematch001_in_chars_last;
  Kernel_inst_rematch001_in_chars                       <= rematch001_in_chars;
  Kernel_inst_rematch001_in_chars_count                 <= rematch001_in_chars_count;

  Kernel_inst_rematch001_in_unl_valid                   <= rematch001_in_unl_valid;
  rematch001_in_unl_ready                               <= Kernel_inst_rematch001_in_unl_ready;
  Kernel_inst_rematch001_in_unl_tag                     <= rematch001_in_unl_tag;

  Kernel_inst_rematch002_in_valid                       <= rematch002_in_valid;
  rematch002_in_ready                                   <= Kernel_inst_rematch002_in_ready;
  Kernel_inst_rematch002_in_dvalid                      <= rematch002_in_dvalid;
  Kernel_inst_rematch002_in_last                        <= rematch002_in_last;
  Kernel_inst_rematch002_in_length                      <= rematch002_in_length;
  Kernel_inst_rematch002_in_count                       <= rematch002_in_count;
  Kernel_inst_rematch002_in_chars_valid                 <= rematch002_in_chars_valid;
  rematch002_in_chars_ready                             <= Kernel_inst_rematch002_in_chars_ready;
  Kernel_inst_rematch002_in_chars_dvalid                <= rematch002_in_chars_dvalid;
  Kernel_inst_rematch002_in_chars_last                  <= rematch002_in_chars_last;
  Kernel_inst_rematch002_in_chars                       <= rematch002_in_chars;
  Kernel_inst_rematch002_in_chars_count                 <= rematch002_in_chars_count;

  Kernel_inst_rematch002_in_unl_valid                   <= rematch002_in_unl_valid;
  rematch002_in_unl_ready                               <= Kernel_inst_rematch002_in_unl_ready;
  Kernel_inst_rematch002_in_unl_tag                     <= rematch002_in_unl_tag;

  Kernel_inst_rematch003_in_valid                       <= rematch003_in_valid;
  rematch003_in_ready                                   <= Kernel_inst_rematch003_in_ready;
  Kernel_inst_rematch003_in_dvalid                      <= rematch003_in_dvalid;
  Kernel_inst_rematch003_in_last                        <= rematch003_in_last;
  Kernel_inst_rematch003_in_length                      <= rematch003_in_length;
  Kernel_inst_rematch003_in_count                       <= rematch003_in_count;
  Kernel_inst_rematch003_in_chars_valid                 <= rematch003_in_chars_valid;
  rematch003_in_chars_ready                             <= Kernel_inst_rematch003_in_chars_ready;
  Kernel_inst_rematch003_in_chars_dvalid                <= rematch003_in_chars_dvalid;
  Kernel_inst_rematch003_in_chars_last                  <= rematch003_in_chars_last;
  Kernel_inst_rematch003_in_chars                       <= rematch003_in_chars;
  Kernel_inst_rematch003_in_chars_count                 <= rematch003_in_chars_count;

  Kernel_inst_rematch003_in_unl_valid                   <= rematch003_in_unl_valid;
  rematch003_in_unl_ready                               <= Kernel_inst_rematch003_in_unl_ready;
  Kernel_inst_rematch003_in_unl_tag                     <= rematch003_in_unl_tag;

  Kernel_inst_rematch004_in_valid                       <= rematch004_in_valid;
  rematch004_in_ready                                   <= Kernel_inst_rematch004_in_ready;
  Kernel_inst_rematch004_in_dvalid                      <= rematch004_in_dvalid;
  Kernel_inst_rematch004_in_last                        <= rematch004_in_last;
  Kernel_inst_rematch004_in_length                      <= rematch004_in_length;
  Kernel_inst_rematch004_in_count                       <= rematch004_in_count;
  Kernel_inst_rematch004_in_chars_valid                 <= rematch004_in_chars_valid;
  rematch004_in_chars_ready                             <= Kernel_inst_rematch004_in_chars_ready;
  Kernel_inst_rematch004_in_chars_dvalid                <= rematch004_in_chars_dvalid;
  Kernel_inst_rematch004_in_chars_last                  <= rematch004_in_chars_last;
  Kernel_inst_rematch004_in_chars                       <= rematch004_in_chars;
  Kernel_inst_rematch004_in_chars_count                 <= rematch004_in_chars_count;

  Kernel_inst_rematch004_in_unl_valid                   <= rematch004_in_unl_valid;
  rematch004_in_unl_ready                               <= Kernel_inst_rematch004_in_unl_ready;
  Kernel_inst_rematch004_in_unl_tag                     <= rematch004_in_unl_tag;

  Kernel_inst_rematch005_in_valid                       <= rematch005_in_valid;
  rematch005_in_ready                                   <= Kernel_inst_rematch005_in_ready;
  Kernel_inst_rematch005_in_dvalid                      <= rematch005_in_dvalid;
  Kernel_inst_rematch005_in_last                        <= rematch005_in_last;
  Kernel_inst_rematch005_in_length                      <= rematch005_in_length;
  Kernel_inst_rematch005_in_count                       <= rematch005_in_count;
  Kernel_inst_rematch005_in_chars_valid                 <= rematch005_in_chars_valid;
  rematch005_in_chars_ready                             <= Kernel_inst_rematch005_in_chars_ready;
  Kernel_inst_rematch005_in_chars_dvalid                <= rematch005_in_chars_dvalid;
  Kernel_inst_rematch005_in_chars_last                  <= rematch005_in_chars_last;
  Kernel_inst_rematch005_in_chars                       <= rematch005_in_chars;
  Kernel_inst_rematch005_in_chars_count                 <= rematch005_in_chars_count;

  Kernel_inst_rematch005_in_unl_valid                   <= rematch005_in_unl_valid;
  rematch005_in_unl_ready                               <= Kernel_inst_rematch005_in_unl_ready;
  Kernel_inst_rematch005_in_unl_tag                     <= rematch005_in_unl_tag;

  Kernel_inst_rematch006_in_valid                       <= rematch006_in_valid;
  rematch006_in_ready                                   <= Kernel_inst_rematch006_in_ready;
  Kernel_inst_rematch006_in_dvalid                      <= rematch006_in_dvalid;
  Kernel_inst_rematch006_in_last                        <= rematch006_in_last;
  Kernel_inst_rematch006_in_length                      <= rematch006_in_length;
  Kernel_inst_rematch006_in_count                       <= rematch006_in_count;
  Kernel_inst_rematch006_in_chars_valid                 <= rematch006_in_chars_valid;
  rematch006_in_chars_ready                             <= Kernel_inst_rematch006_in_chars_ready;
  Kernel_inst_rematch006_in_chars_dvalid                <= rematch006_in_chars_dvalid;
  Kernel_inst_rematch006_in_chars_last                  <= rematch006_in_chars_last;
  Kernel_inst_rematch006_in_chars                       <= rematch006_in_chars;
  Kernel_inst_rematch006_in_chars_count                 <= rematch006_in_chars_count;

  Kernel_inst_rematch006_in_unl_valid                   <= rematch006_in_unl_valid;
  rematch006_in_unl_ready                               <= Kernel_inst_rematch006_in_unl_ready;
  Kernel_inst_rematch006_in_unl_tag                     <= rematch006_in_unl_tag;

  Kernel_inst_rematch007_in_valid                       <= rematch007_in_valid;
  rematch007_in_ready                                   <= Kernel_inst_rematch007_in_ready;
  Kernel_inst_rematch007_in_dvalid                      <= rematch007_in_dvalid;
  Kernel_inst_rematch007_in_last                        <= rematch007_in_last;
  Kernel_inst_rematch007_in_length                      <= rematch007_in_length;
  Kernel_inst_rematch007_in_count                       <= rematch007_in_count;
  Kernel_inst_rematch007_in_chars_valid                 <= rematch007_in_chars_valid;
  rematch007_in_chars_ready                             <= Kernel_inst_rematch007_in_chars_ready;
  Kernel_inst_rematch007_in_chars_dvalid                <= rematch007_in_chars_dvalid;
  Kernel_inst_rematch007_in_chars_last                  <= rematch007_in_chars_last;
  Kernel_inst_rematch007_in_chars                       <= rematch007_in_chars;
  Kernel_inst_rematch007_in_chars_count                 <= rematch007_in_chars_count;

  Kernel_inst_rematch007_in_unl_valid                   <= rematch007_in_unl_valid;
  rematch007_in_unl_ready                               <= Kernel_inst_rematch007_in_unl_ready;
  Kernel_inst_rematch007_in_unl_tag                     <= rematch007_in_unl_tag;

  Kernel_inst_rematch008_in_valid                       <= rematch008_in_valid;
  rematch008_in_ready                                   <= Kernel_inst_rematch008_in_ready;
  Kernel_inst_rematch008_in_dvalid                      <= rematch008_in_dvalid;
  Kernel_inst_rematch008_in_last                        <= rematch008_in_last;
  Kernel_inst_rematch008_in_length                      <= rematch008_in_length;
  Kernel_inst_rematch008_in_count                       <= rematch008_in_count;
  Kernel_inst_rematch008_in_chars_valid                 <= rematch008_in_chars_valid;
  rematch008_in_chars_ready                             <= Kernel_inst_rematch008_in_chars_ready;
  Kernel_inst_rematch008_in_chars_dvalid                <= rematch008_in_chars_dvalid;
  Kernel_inst_rematch008_in_chars_last                  <= rematch008_in_chars_last;
  Kernel_inst_rematch008_in_chars                       <= rematch008_in_chars;
  Kernel_inst_rematch008_in_chars_count                 <= rematch008_in_chars_count;

  Kernel_inst_rematch008_in_unl_valid                   <= rematch008_in_unl_valid;
  rematch008_in_unl_ready                               <= Kernel_inst_rematch008_in_unl_ready;
  Kernel_inst_rematch008_in_unl_tag                     <= rematch008_in_unl_tag;

  Kernel_inst_rematch009_in_valid                       <= rematch009_in_valid;
  rematch009_in_ready                                   <= Kernel_inst_rematch009_in_ready;
  Kernel_inst_rematch009_in_dvalid                      <= rematch009_in_dvalid;
  Kernel_inst_rematch009_in_last                        <= rematch009_in_last;
  Kernel_inst_rematch009_in_length                      <= rematch009_in_length;
  Kernel_inst_rematch009_in_count                       <= rematch009_in_count;
  Kernel_inst_rematch009_in_chars_valid                 <= rematch009_in_chars_valid;
  rematch009_in_chars_ready                             <= Kernel_inst_rematch009_in_chars_ready;
  Kernel_inst_rematch009_in_chars_dvalid                <= rematch009_in_chars_dvalid;
  Kernel_inst_rematch009_in_chars_last                  <= rematch009_in_chars_last;
  Kernel_inst_rematch009_in_chars                       <= rematch009_in_chars;
  Kernel_inst_rematch009_in_chars_count                 <= rematch009_in_chars_count;

  Kernel_inst_rematch009_in_unl_valid                   <= rematch009_in_unl_valid;
  rematch009_in_unl_ready                               <= Kernel_inst_rematch009_in_unl_ready;
  Kernel_inst_rematch009_in_unl_tag                     <= rematch009_in_unl_tag;

  Kernel_inst_rematch010_in_valid                       <= rematch010_in_valid;
  rematch010_in_ready                                   <= Kernel_inst_rematch010_in_ready;
  Kernel_inst_rematch010_in_dvalid                      <= rematch010_in_dvalid;
  Kernel_inst_rematch010_in_last                        <= rematch010_in_last;
  Kernel_inst_rematch010_in_length                      <= rematch010_in_length;
  Kernel_inst_rematch010_in_count                       <= rematch010_in_count;
  Kernel_inst_rematch010_in_chars_valid                 <= rematch010_in_chars_valid;
  rematch010_in_chars_ready                             <= Kernel_inst_rematch010_in_chars_ready;
  Kernel_inst_rematch010_in_chars_dvalid                <= rematch010_in_chars_dvalid;
  Kernel_inst_rematch010_in_chars_last                  <= rematch010_in_chars_last;
  Kernel_inst_rematch010_in_chars                       <= rematch010_in_chars;
  Kernel_inst_rematch010_in_chars_count                 <= rematch010_in_chars_count;

  Kernel_inst_rematch010_in_unl_valid                   <= rematch010_in_unl_valid;
  rematch010_in_unl_ready                               <= Kernel_inst_rematch010_in_unl_ready;
  Kernel_inst_rematch010_in_unl_tag                     <= rematch010_in_unl_tag;

  Kernel_inst_rematch011_in_valid                       <= rematch011_in_valid;
  rematch011_in_ready                                   <= Kernel_inst_rematch011_in_ready;
  Kernel_inst_rematch011_in_dvalid                      <= rematch011_in_dvalid;
  Kernel_inst_rematch011_in_last                        <= rematch011_in_last;
  Kernel_inst_rematch011_in_length                      <= rematch011_in_length;
  Kernel_inst_rematch011_in_count                       <= rematch011_in_count;
  Kernel_inst_rematch011_in_chars_valid                 <= rematch011_in_chars_valid;
  rematch011_in_chars_ready                             <= Kernel_inst_rematch011_in_chars_ready;
  Kernel_inst_rematch011_in_chars_dvalid                <= rematch011_in_chars_dvalid;
  Kernel_inst_rematch011_in_chars_last                  <= rematch011_in_chars_last;
  Kernel_inst_rematch011_in_chars                       <= rematch011_in_chars;
  Kernel_inst_rematch011_in_chars_count                 <= rematch011_in_chars_count;

  Kernel_inst_rematch011_in_unl_valid                   <= rematch011_in_unl_valid;
  rematch011_in_unl_ready                               <= Kernel_inst_rematch011_in_unl_ready;
  Kernel_inst_rematch011_in_unl_tag                     <= rematch011_in_unl_tag;

  Kernel_inst_rematch012_in_valid                       <= rematch012_in_valid;
  rematch012_in_ready                                   <= Kernel_inst_rematch012_in_ready;
  Kernel_inst_rematch012_in_dvalid                      <= rematch012_in_dvalid;
  Kernel_inst_rematch012_in_last                        <= rematch012_in_last;
  Kernel_inst_rematch012_in_length                      <= rematch012_in_length;
  Kernel_inst_rematch012_in_count                       <= rematch012_in_count;
  Kernel_inst_rematch012_in_chars_valid                 <= rematch012_in_chars_valid;
  rematch012_in_chars_ready                             <= Kernel_inst_rematch012_in_chars_ready;
  Kernel_inst_rematch012_in_chars_dvalid                <= rematch012_in_chars_dvalid;
  Kernel_inst_rematch012_in_chars_last                  <= rematch012_in_chars_last;
  Kernel_inst_rematch012_in_chars                       <= rematch012_in_chars;
  Kernel_inst_rematch012_in_chars_count                 <= rematch012_in_chars_count;

  Kernel_inst_rematch012_in_unl_valid                   <= rematch012_in_unl_valid;
  rematch012_in_unl_ready                               <= Kernel_inst_rematch012_in_unl_ready;
  Kernel_inst_rematch012_in_unl_tag                     <= rematch012_in_unl_tag;

  Kernel_inst_rematch013_in_valid                       <= rematch013_in_valid;
  rematch013_in_ready                                   <= Kernel_inst_rematch013_in_ready;
  Kernel_inst_rematch013_in_dvalid                      <= rematch013_in_dvalid;
  Kernel_inst_rematch013_in_last                        <= rematch013_in_last;
  Kernel_inst_rematch013_in_length                      <= rematch013_in_length;
  Kernel_inst_rematch013_in_count                       <= rematch013_in_count;
  Kernel_inst_rematch013_in_chars_valid                 <= rematch013_in_chars_valid;
  rematch013_in_chars_ready                             <= Kernel_inst_rematch013_in_chars_ready;
  Kernel_inst_rematch013_in_chars_dvalid                <= rematch013_in_chars_dvalid;
  Kernel_inst_rematch013_in_chars_last                  <= rematch013_in_chars_last;
  Kernel_inst_rematch013_in_chars                       <= rematch013_in_chars;
  Kernel_inst_rematch013_in_chars_count                 <= rematch013_in_chars_count;

  Kernel_inst_rematch013_in_unl_valid                   <= rematch013_in_unl_valid;
  rematch013_in_unl_ready                               <= Kernel_inst_rematch013_in_unl_ready;
  Kernel_inst_rematch013_in_unl_tag                     <= rematch013_in_unl_tag;

  Kernel_inst_rematch014_in_valid                       <= rematch014_in_valid;
  rematch014_in_ready                                   <= Kernel_inst_rematch014_in_ready;
  Kernel_inst_rematch014_in_dvalid                      <= rematch014_in_dvalid;
  Kernel_inst_rematch014_in_last                        <= rematch014_in_last;
  Kernel_inst_rematch014_in_length                      <= rematch014_in_length;
  Kernel_inst_rematch014_in_count                       <= rematch014_in_count;
  Kernel_inst_rematch014_in_chars_valid                 <= rematch014_in_chars_valid;
  rematch014_in_chars_ready                             <= Kernel_inst_rematch014_in_chars_ready;
  Kernel_inst_rematch014_in_chars_dvalid                <= rematch014_in_chars_dvalid;
  Kernel_inst_rematch014_in_chars_last                  <= rematch014_in_chars_last;
  Kernel_inst_rematch014_in_chars                       <= rematch014_in_chars;
  Kernel_inst_rematch014_in_chars_count                 <= rematch014_in_chars_count;

  Kernel_inst_rematch014_in_unl_valid                   <= rematch014_in_unl_valid;
  rematch014_in_unl_ready                               <= Kernel_inst_rematch014_in_unl_ready;
  Kernel_inst_rematch014_in_unl_tag                     <= rematch014_in_unl_tag;

  Kernel_inst_rematch015_in_valid                       <= rematch015_in_valid;
  rematch015_in_ready                                   <= Kernel_inst_rematch015_in_ready;
  Kernel_inst_rematch015_in_dvalid                      <= rematch015_in_dvalid;
  Kernel_inst_rematch015_in_last                        <= rematch015_in_last;
  Kernel_inst_rematch015_in_length                      <= rematch015_in_length;
  Kernel_inst_rematch015_in_count                       <= rematch015_in_count;
  Kernel_inst_rematch015_in_chars_valid                 <= rematch015_in_chars_valid;
  rematch015_in_chars_ready                             <= Kernel_inst_rematch015_in_chars_ready;
  Kernel_inst_rematch015_in_chars_dvalid                <= rematch015_in_chars_dvalid;
  Kernel_inst_rematch015_in_chars_last                  <= rematch015_in_chars_last;
  Kernel_inst_rematch015_in_chars                       <= rematch015_in_chars;
  Kernel_inst_rematch015_in_chars_count                 <= rematch015_in_chars_count;

  Kernel_inst_rematch015_in_unl_valid                   <= rematch015_in_unl_valid;
  rematch015_in_unl_ready                               <= Kernel_inst_rematch015_in_unl_ready;
  Kernel_inst_rematch015_in_unl_tag                     <= rematch015_in_unl_tag;

  Kernel_inst_rematch000_taxi_out_unl_valid             <= rematch000_taxi_out_unl_valid;
  rematch000_taxi_out_unl_ready                         <= Kernel_inst_rematch000_taxi_out_unl_ready;
  Kernel_inst_rematch000_taxi_out_unl_tag               <= rematch000_taxi_out_unl_tag;

  Kernel_inst_rematch001_taxi_out_unl_valid             <= rematch001_taxi_out_unl_valid;
  rematch001_taxi_out_unl_ready                         <= Kernel_inst_rematch001_taxi_out_unl_ready;
  Kernel_inst_rematch001_taxi_out_unl_tag               <= rematch001_taxi_out_unl_tag;

  Kernel_inst_rematch002_taxi_out_unl_valid             <= rematch002_taxi_out_unl_valid;
  rematch002_taxi_out_unl_ready                         <= Kernel_inst_rematch002_taxi_out_unl_ready;
  Kernel_inst_rematch002_taxi_out_unl_tag               <= rematch002_taxi_out_unl_tag;

  Kernel_inst_rematch003_taxi_out_unl_valid             <= rematch003_taxi_out_unl_valid;
  rematch003_taxi_out_unl_ready                         <= Kernel_inst_rematch003_taxi_out_unl_ready;
  Kernel_inst_rematch003_taxi_out_unl_tag               <= rematch003_taxi_out_unl_tag;

  Kernel_inst_rematch004_taxi_out_unl_valid             <= rematch004_taxi_out_unl_valid;
  rematch004_taxi_out_unl_ready                         <= Kernel_inst_rematch004_taxi_out_unl_ready;
  Kernel_inst_rematch004_taxi_out_unl_tag               <= rematch004_taxi_out_unl_tag;

  Kernel_inst_rematch005_taxi_out_unl_valid             <= rematch005_taxi_out_unl_valid;
  rematch005_taxi_out_unl_ready                         <= Kernel_inst_rematch005_taxi_out_unl_ready;
  Kernel_inst_rematch005_taxi_out_unl_tag               <= rematch005_taxi_out_unl_tag;

  Kernel_inst_rematch006_taxi_out_unl_valid             <= rematch006_taxi_out_unl_valid;
  rematch006_taxi_out_unl_ready                         <= Kernel_inst_rematch006_taxi_out_unl_ready;
  Kernel_inst_rematch006_taxi_out_unl_tag               <= rematch006_taxi_out_unl_tag;

  Kernel_inst_rematch007_taxi_out_unl_valid             <= rematch007_taxi_out_unl_valid;
  rematch007_taxi_out_unl_ready                         <= Kernel_inst_rematch007_taxi_out_unl_ready;
  Kernel_inst_rematch007_taxi_out_unl_tag               <= rematch007_taxi_out_unl_tag;

  Kernel_inst_rematch008_taxi_out_unl_valid             <= rematch008_taxi_out_unl_valid;
  rematch008_taxi_out_unl_ready                         <= Kernel_inst_rematch008_taxi_out_unl_ready;
  Kernel_inst_rematch008_taxi_out_unl_tag               <= rematch008_taxi_out_unl_tag;

  Kernel_inst_rematch009_taxi_out_unl_valid             <= rematch009_taxi_out_unl_valid;
  rematch009_taxi_out_unl_ready                         <= Kernel_inst_rematch009_taxi_out_unl_ready;
  Kernel_inst_rematch009_taxi_out_unl_tag               <= rematch009_taxi_out_unl_tag;

  Kernel_inst_rematch010_taxi_out_unl_valid             <= rematch010_taxi_out_unl_valid;
  rematch010_taxi_out_unl_ready                         <= Kernel_inst_rematch010_taxi_out_unl_ready;
  Kernel_inst_rematch010_taxi_out_unl_tag               <= rematch010_taxi_out_unl_tag;

  Kernel_inst_rematch011_taxi_out_unl_valid             <= rematch011_taxi_out_unl_valid;
  rematch011_taxi_out_unl_ready                         <= Kernel_inst_rematch011_taxi_out_unl_ready;
  Kernel_inst_rematch011_taxi_out_unl_tag               <= rematch011_taxi_out_unl_tag;

  Kernel_inst_rematch012_taxi_out_unl_valid             <= rematch012_taxi_out_unl_valid;
  rematch012_taxi_out_unl_ready                         <= Kernel_inst_rematch012_taxi_out_unl_ready;
  Kernel_inst_rematch012_taxi_out_unl_tag               <= rematch012_taxi_out_unl_tag;

  Kernel_inst_rematch013_taxi_out_unl_valid             <= rematch013_taxi_out_unl_valid;
  rematch013_taxi_out_unl_ready                         <= Kernel_inst_rematch013_taxi_out_unl_ready;
  Kernel_inst_rematch013_taxi_out_unl_tag               <= rematch013_taxi_out_unl_tag;

  Kernel_inst_rematch014_taxi_out_unl_valid             <= rematch014_taxi_out_unl_valid;
  rematch014_taxi_out_unl_ready                         <= Kernel_inst_rematch014_taxi_out_unl_ready;
  Kernel_inst_rematch014_taxi_out_unl_tag               <= rematch014_taxi_out_unl_tag;

  Kernel_inst_rematch015_taxi_out_unl_valid             <= rematch015_taxi_out_unl_valid;
  rematch015_taxi_out_unl_ready                         <= Kernel_inst_rematch015_taxi_out_unl_ready;
  Kernel_inst_rematch015_taxi_out_unl_tag               <= rematch015_taxi_out_unl_tag;

  Kernel_inst_start                                     <= mmio_inst_f_start_data;
  Kernel_inst_stop                                      <= mmio_inst_f_stop_data;
  Kernel_inst_reset                                     <= mmio_inst_f_reset_data;
  Kernel_inst_rematch000_firstidx                       <= mmio_inst_f_rematch000_firstidx_data;
  Kernel_inst_rematch000_lastidx                        <= mmio_inst_f_rematch000_lastidx_data;
  Kernel_inst_rematch001_firstidx                       <= mmio_inst_f_rematch001_firstidx_data;
  Kernel_inst_rematch001_lastidx                        <= mmio_inst_f_rematch001_lastidx_data;
  Kernel_inst_rematch002_firstidx                       <= mmio_inst_f_rematch002_firstidx_data;
  Kernel_inst_rematch002_lastidx                        <= mmio_inst_f_rematch002_lastidx_data;
  Kernel_inst_rematch003_firstidx                       <= mmio_inst_f_rematch003_firstidx_data;
  Kernel_inst_rematch003_lastidx                        <= mmio_inst_f_rematch003_lastidx_data;
  Kernel_inst_rematch004_firstidx                       <= mmio_inst_f_rematch004_firstidx_data;
  Kernel_inst_rematch004_lastidx                        <= mmio_inst_f_rematch004_lastidx_data;
  Kernel_inst_rematch005_firstidx                       <= mmio_inst_f_rematch005_firstidx_data;
  Kernel_inst_rematch005_lastidx                        <= mmio_inst_f_rematch005_lastidx_data;
  Kernel_inst_rematch006_firstidx                       <= mmio_inst_f_rematch006_firstidx_data;
  Kernel_inst_rematch006_lastidx                        <= mmio_inst_f_rematch006_lastidx_data;
  Kernel_inst_rematch007_firstidx                       <= mmio_inst_f_rematch007_firstidx_data;
  Kernel_inst_rematch007_lastidx                        <= mmio_inst_f_rematch007_lastidx_data;
  Kernel_inst_rematch008_firstidx                       <= mmio_inst_f_rematch008_firstidx_data;
  Kernel_inst_rematch008_lastidx                        <= mmio_inst_f_rematch008_lastidx_data;
  Kernel_inst_rematch009_firstidx                       <= mmio_inst_f_rematch009_firstidx_data;
  Kernel_inst_rematch009_lastidx                        <= mmio_inst_f_rematch009_lastidx_data;
  Kernel_inst_rematch010_firstidx                       <= mmio_inst_f_rematch010_firstidx_data;
  Kernel_inst_rematch010_lastidx                        <= mmio_inst_f_rematch010_lastidx_data;
  Kernel_inst_rematch011_firstidx                       <= mmio_inst_f_rematch011_firstidx_data;
  Kernel_inst_rematch011_lastidx                        <= mmio_inst_f_rematch011_lastidx_data;
  Kernel_inst_rematch012_firstidx                       <= mmio_inst_f_rematch012_firstidx_data;
  Kernel_inst_rematch012_lastidx                        <= mmio_inst_f_rematch012_lastidx_data;
  Kernel_inst_rematch013_firstidx                       <= mmio_inst_f_rematch013_firstidx_data;
  Kernel_inst_rematch013_lastidx                        <= mmio_inst_f_rematch013_lastidx_data;
  Kernel_inst_rematch014_firstidx                       <= mmio_inst_f_rematch014_firstidx_data;
  Kernel_inst_rematch014_lastidx                        <= mmio_inst_f_rematch014_lastidx_data;
  Kernel_inst_rematch015_firstidx                       <= mmio_inst_f_rematch015_firstidx_data;
  Kernel_inst_rematch015_lastidx                        <= mmio_inst_f_rematch015_lastidx_data;
  Kernel_inst_rematch000_taxi_firstidx                  <= mmio_inst_f_rematch000_taxi_firstidx_data;
  Kernel_inst_rematch000_taxi_lastidx                   <= mmio_inst_f_rematch000_taxi_lastidx_data;
  Kernel_inst_rematch001_taxi_firstidx                  <= mmio_inst_f_rematch001_taxi_firstidx_data;
  Kernel_inst_rematch001_taxi_lastidx                   <= mmio_inst_f_rematch001_taxi_lastidx_data;
  Kernel_inst_rematch002_taxi_firstidx                  <= mmio_inst_f_rematch002_taxi_firstidx_data;
  Kernel_inst_rematch002_taxi_lastidx                   <= mmio_inst_f_rematch002_taxi_lastidx_data;
  Kernel_inst_rematch003_taxi_firstidx                  <= mmio_inst_f_rematch003_taxi_firstidx_data;
  Kernel_inst_rematch003_taxi_lastidx                   <= mmio_inst_f_rematch003_taxi_lastidx_data;
  Kernel_inst_rematch004_taxi_firstidx                  <= mmio_inst_f_rematch004_taxi_firstidx_data;
  Kernel_inst_rematch004_taxi_lastidx                   <= mmio_inst_f_rematch004_taxi_lastidx_data;
  Kernel_inst_rematch005_taxi_firstidx                  <= mmio_inst_f_rematch005_taxi_firstidx_data;
  Kernel_inst_rematch005_taxi_lastidx                   <= mmio_inst_f_rematch005_taxi_lastidx_data;
  Kernel_inst_rematch006_taxi_firstidx                  <= mmio_inst_f_rematch006_taxi_firstidx_data;
  Kernel_inst_rematch006_taxi_lastidx                   <= mmio_inst_f_rematch006_taxi_lastidx_data;
  Kernel_inst_rematch007_taxi_firstidx                  <= mmio_inst_f_rematch007_taxi_firstidx_data;
  Kernel_inst_rematch007_taxi_lastidx                   <= mmio_inst_f_rematch007_taxi_lastidx_data;
  Kernel_inst_rematch008_taxi_firstidx                  <= mmio_inst_f_rematch008_taxi_firstidx_data;
  Kernel_inst_rematch008_taxi_lastidx                   <= mmio_inst_f_rematch008_taxi_lastidx_data;
  Kernel_inst_rematch009_taxi_firstidx                  <= mmio_inst_f_rematch009_taxi_firstidx_data;
  Kernel_inst_rematch009_taxi_lastidx                   <= mmio_inst_f_rematch009_taxi_lastidx_data;
  Kernel_inst_rematch010_taxi_firstidx                  <= mmio_inst_f_rematch010_taxi_firstidx_data;
  Kernel_inst_rematch010_taxi_lastidx                   <= mmio_inst_f_rematch010_taxi_lastidx_data;
  Kernel_inst_rematch011_taxi_firstidx                  <= mmio_inst_f_rematch011_taxi_firstidx_data;
  Kernel_inst_rematch011_taxi_lastidx                   <= mmio_inst_f_rematch011_taxi_lastidx_data;
  Kernel_inst_rematch012_taxi_firstidx                  <= mmio_inst_f_rematch012_taxi_firstidx_data;
  Kernel_inst_rematch012_taxi_lastidx                   <= mmio_inst_f_rematch012_taxi_lastidx_data;
  Kernel_inst_rematch013_taxi_firstidx                  <= mmio_inst_f_rematch013_taxi_firstidx_data;
  Kernel_inst_rematch013_taxi_lastidx                   <= mmio_inst_f_rematch013_taxi_lastidx_data;
  Kernel_inst_rematch014_taxi_firstidx                  <= mmio_inst_f_rematch014_taxi_firstidx_data;
  Kernel_inst_rematch014_taxi_lastidx                   <= mmio_inst_f_rematch014_taxi_lastidx_data;
  Kernel_inst_rematch015_taxi_firstidx                  <= mmio_inst_f_rematch015_taxi_firstidx_data;
  Kernel_inst_rematch015_taxi_lastidx                   <= mmio_inst_f_rematch015_taxi_lastidx_data;
  mmio_inst_f_idle_write_data                           <= Kernel_inst_idle;
  mmio_inst_f_busy_write_data                           <= Kernel_inst_busy;
  mmio_inst_f_done_write_data                           <= Kernel_inst_done;
  mmio_inst_f_result_write_data                         <= Kernel_inst_result;
  mmio_inst_f_rematch000_taxi_count_write_data          <= Kernel_inst_rematch000_taxi_count;
  mmio_inst_f_rematch000_errors_write_data              <= Kernel_inst_rematch000_errors;
  mmio_inst_f_rematch001_taxi_count_write_data          <= Kernel_inst_rematch001_taxi_count;
  mmio_inst_f_rematch001_errors_write_data              <= Kernel_inst_rematch001_errors;
  mmio_inst_f_rematch002_taxi_count_write_data          <= Kernel_inst_rematch002_taxi_count;
  mmio_inst_f_rematch002_errors_write_data              <= Kernel_inst_rematch002_errors;
  mmio_inst_f_rematch003_taxi_count_write_data          <= Kernel_inst_rematch003_taxi_count;
  mmio_inst_f_rematch003_errors_write_data              <= Kernel_inst_rematch003_errors;
  mmio_inst_f_rematch004_taxi_count_write_data          <= Kernel_inst_rematch004_taxi_count;
  mmio_inst_f_rematch004_errors_write_data              <= Kernel_inst_rematch004_errors;
  mmio_inst_f_rematch005_taxi_count_write_data          <= Kernel_inst_rematch005_taxi_count;
  mmio_inst_f_rematch005_errors_write_data              <= Kernel_inst_rematch005_errors;
  mmio_inst_f_rematch006_taxi_count_write_data          <= Kernel_inst_rematch006_taxi_count;
  mmio_inst_f_rematch006_errors_write_data              <= Kernel_inst_rematch006_errors;
  mmio_inst_f_rematch007_taxi_count_write_data          <= Kernel_inst_rematch007_taxi_count;
  mmio_inst_f_rematch007_errors_write_data              <= Kernel_inst_rematch007_errors;
  mmio_inst_f_rematch008_taxi_count_write_data          <= Kernel_inst_rematch008_taxi_count;
  mmio_inst_f_rematch008_errors_write_data              <= Kernel_inst_rematch008_errors;
  mmio_inst_f_rematch009_taxi_count_write_data          <= Kernel_inst_rematch009_taxi_count;
  mmio_inst_f_rematch009_errors_write_data              <= Kernel_inst_rematch009_errors;
  mmio_inst_f_rematch010_taxi_count_write_data          <= Kernel_inst_rematch010_taxi_count;
  mmio_inst_f_rematch010_errors_write_data              <= Kernel_inst_rematch010_errors;
  mmio_inst_f_rematch011_taxi_count_write_data          <= Kernel_inst_rematch011_taxi_count;
  mmio_inst_f_rematch011_errors_write_data              <= Kernel_inst_rematch011_errors;
  mmio_inst_f_rematch012_taxi_count_write_data          <= Kernel_inst_rematch012_taxi_count;
  mmio_inst_f_rematch012_errors_write_data              <= Kernel_inst_rematch012_errors;
  mmio_inst_f_rematch013_taxi_count_write_data          <= Kernel_inst_rematch013_taxi_count;
  mmio_inst_f_rematch013_errors_write_data              <= Kernel_inst_rematch013_errors;
  mmio_inst_f_rematch014_taxi_count_write_data          <= Kernel_inst_rematch014_taxi_count;
  mmio_inst_f_rematch014_errors_write_data              <= Kernel_inst_rematch014_errors;
  mmio_inst_f_rematch015_taxi_count_write_data          <= Kernel_inst_rematch015_taxi_count;
  mmio_inst_f_rematch015_errors_write_data              <= Kernel_inst_rematch015_errors;
  mmio_inst_mmio_awvalid                                <= mmio_awvalid;
  mmio_awready                                          <= mmio_inst_mmio_awready;
  mmio_inst_mmio_awaddr                                 <= mmio_awaddr;
  mmio_inst_mmio_wvalid                                 <= mmio_wvalid;
  mmio_wready                                           <= mmio_inst_mmio_wready;
  mmio_inst_mmio_wdata                                  <= mmio_wdata;
  mmio_inst_mmio_wstrb                                  <= mmio_wstrb;
  mmio_bvalid                                           <= mmio_inst_mmio_bvalid;
  mmio_inst_mmio_bready                                 <= mmio_bready;
  mmio_bresp                                            <= mmio_inst_mmio_bresp;
  mmio_inst_mmio_arvalid                                <= mmio_arvalid;
  mmio_arready                                          <= mmio_inst_mmio_arready;
  mmio_inst_mmio_araddr                                 <= mmio_araddr;
  mmio_rvalid                                           <= mmio_inst_mmio_rvalid;
  mmio_inst_mmio_rready                                 <= mmio_rready;
  mmio_rdata                                            <= mmio_inst_mmio_rdata;
  mmio_rresp                                            <= mmio_inst_mmio_rresp;

  rematch000_in_cmd_accm_inst_kernel_cmd_valid          <= Kernel_inst_rematch000_in_cmd_valid;
  Kernel_inst_rematch000_in_cmd_ready                   <= rematch000_in_cmd_accm_inst_kernel_cmd_ready;
  rematch000_in_cmd_accm_inst_kernel_cmd_firstIdx       <= Kernel_inst_rematch000_in_cmd_firstIdx;
  rematch000_in_cmd_accm_inst_kernel_cmd_lastIdx        <= Kernel_inst_rematch000_in_cmd_lastIdx;
  rematch000_in_cmd_accm_inst_kernel_cmd_tag            <= Kernel_inst_rematch000_in_cmd_tag;

  rematch001_in_cmd_accm_inst_kernel_cmd_valid          <= Kernel_inst_rematch001_in_cmd_valid;
  Kernel_inst_rematch001_in_cmd_ready                   <= rematch001_in_cmd_accm_inst_kernel_cmd_ready;
  rematch001_in_cmd_accm_inst_kernel_cmd_firstIdx       <= Kernel_inst_rematch001_in_cmd_firstIdx;
  rematch001_in_cmd_accm_inst_kernel_cmd_lastIdx        <= Kernel_inst_rematch001_in_cmd_lastIdx;
  rematch001_in_cmd_accm_inst_kernel_cmd_tag            <= Kernel_inst_rematch001_in_cmd_tag;

  rematch002_in_cmd_accm_inst_kernel_cmd_valid          <= Kernel_inst_rematch002_in_cmd_valid;
  Kernel_inst_rematch002_in_cmd_ready                   <= rematch002_in_cmd_accm_inst_kernel_cmd_ready;
  rematch002_in_cmd_accm_inst_kernel_cmd_firstIdx       <= Kernel_inst_rematch002_in_cmd_firstIdx;
  rematch002_in_cmd_accm_inst_kernel_cmd_lastIdx        <= Kernel_inst_rematch002_in_cmd_lastIdx;
  rematch002_in_cmd_accm_inst_kernel_cmd_tag            <= Kernel_inst_rematch002_in_cmd_tag;

  rematch003_in_cmd_accm_inst_kernel_cmd_valid          <= Kernel_inst_rematch003_in_cmd_valid;
  Kernel_inst_rematch003_in_cmd_ready                   <= rematch003_in_cmd_accm_inst_kernel_cmd_ready;
  rematch003_in_cmd_accm_inst_kernel_cmd_firstIdx       <= Kernel_inst_rematch003_in_cmd_firstIdx;
  rematch003_in_cmd_accm_inst_kernel_cmd_lastIdx        <= Kernel_inst_rematch003_in_cmd_lastIdx;
  rematch003_in_cmd_accm_inst_kernel_cmd_tag            <= Kernel_inst_rematch003_in_cmd_tag;

  rematch004_in_cmd_accm_inst_kernel_cmd_valid          <= Kernel_inst_rematch004_in_cmd_valid;
  Kernel_inst_rematch004_in_cmd_ready                   <= rematch004_in_cmd_accm_inst_kernel_cmd_ready;
  rematch004_in_cmd_accm_inst_kernel_cmd_firstIdx       <= Kernel_inst_rematch004_in_cmd_firstIdx;
  rematch004_in_cmd_accm_inst_kernel_cmd_lastIdx        <= Kernel_inst_rematch004_in_cmd_lastIdx;
  rematch004_in_cmd_accm_inst_kernel_cmd_tag            <= Kernel_inst_rematch004_in_cmd_tag;

  rematch005_in_cmd_accm_inst_kernel_cmd_valid          <= Kernel_inst_rematch005_in_cmd_valid;
  Kernel_inst_rematch005_in_cmd_ready                   <= rematch005_in_cmd_accm_inst_kernel_cmd_ready;
  rematch005_in_cmd_accm_inst_kernel_cmd_firstIdx       <= Kernel_inst_rematch005_in_cmd_firstIdx;
  rematch005_in_cmd_accm_inst_kernel_cmd_lastIdx        <= Kernel_inst_rematch005_in_cmd_lastIdx;
  rematch005_in_cmd_accm_inst_kernel_cmd_tag            <= Kernel_inst_rematch005_in_cmd_tag;

  rematch006_in_cmd_accm_inst_kernel_cmd_valid          <= Kernel_inst_rematch006_in_cmd_valid;
  Kernel_inst_rematch006_in_cmd_ready                   <= rematch006_in_cmd_accm_inst_kernel_cmd_ready;
  rematch006_in_cmd_accm_inst_kernel_cmd_firstIdx       <= Kernel_inst_rematch006_in_cmd_firstIdx;
  rematch006_in_cmd_accm_inst_kernel_cmd_lastIdx        <= Kernel_inst_rematch006_in_cmd_lastIdx;
  rematch006_in_cmd_accm_inst_kernel_cmd_tag            <= Kernel_inst_rematch006_in_cmd_tag;

  rematch007_in_cmd_accm_inst_kernel_cmd_valid          <= Kernel_inst_rematch007_in_cmd_valid;
  Kernel_inst_rematch007_in_cmd_ready                   <= rematch007_in_cmd_accm_inst_kernel_cmd_ready;
  rematch007_in_cmd_accm_inst_kernel_cmd_firstIdx       <= Kernel_inst_rematch007_in_cmd_firstIdx;
  rematch007_in_cmd_accm_inst_kernel_cmd_lastIdx        <= Kernel_inst_rematch007_in_cmd_lastIdx;
  rematch007_in_cmd_accm_inst_kernel_cmd_tag            <= Kernel_inst_rematch007_in_cmd_tag;

  rematch008_in_cmd_accm_inst_kernel_cmd_valid          <= Kernel_inst_rematch008_in_cmd_valid;
  Kernel_inst_rematch008_in_cmd_ready                   <= rematch008_in_cmd_accm_inst_kernel_cmd_ready;
  rematch008_in_cmd_accm_inst_kernel_cmd_firstIdx       <= Kernel_inst_rematch008_in_cmd_firstIdx;
  rematch008_in_cmd_accm_inst_kernel_cmd_lastIdx        <= Kernel_inst_rematch008_in_cmd_lastIdx;
  rematch008_in_cmd_accm_inst_kernel_cmd_tag            <= Kernel_inst_rematch008_in_cmd_tag;

  rematch009_in_cmd_accm_inst_kernel_cmd_valid          <= Kernel_inst_rematch009_in_cmd_valid;
  Kernel_inst_rematch009_in_cmd_ready                   <= rematch009_in_cmd_accm_inst_kernel_cmd_ready;
  rematch009_in_cmd_accm_inst_kernel_cmd_firstIdx       <= Kernel_inst_rematch009_in_cmd_firstIdx;
  rematch009_in_cmd_accm_inst_kernel_cmd_lastIdx        <= Kernel_inst_rematch009_in_cmd_lastIdx;
  rematch009_in_cmd_accm_inst_kernel_cmd_tag            <= Kernel_inst_rematch009_in_cmd_tag;

  rematch010_in_cmd_accm_inst_kernel_cmd_valid          <= Kernel_inst_rematch010_in_cmd_valid;
  Kernel_inst_rematch010_in_cmd_ready                   <= rematch010_in_cmd_accm_inst_kernel_cmd_ready;
  rematch010_in_cmd_accm_inst_kernel_cmd_firstIdx       <= Kernel_inst_rematch010_in_cmd_firstIdx;
  rematch010_in_cmd_accm_inst_kernel_cmd_lastIdx        <= Kernel_inst_rematch010_in_cmd_lastIdx;
  rematch010_in_cmd_accm_inst_kernel_cmd_tag            <= Kernel_inst_rematch010_in_cmd_tag;

  rematch011_in_cmd_accm_inst_kernel_cmd_valid          <= Kernel_inst_rematch011_in_cmd_valid;
  Kernel_inst_rematch011_in_cmd_ready                   <= rematch011_in_cmd_accm_inst_kernel_cmd_ready;
  rematch011_in_cmd_accm_inst_kernel_cmd_firstIdx       <= Kernel_inst_rematch011_in_cmd_firstIdx;
  rematch011_in_cmd_accm_inst_kernel_cmd_lastIdx        <= Kernel_inst_rematch011_in_cmd_lastIdx;
  rematch011_in_cmd_accm_inst_kernel_cmd_tag            <= Kernel_inst_rematch011_in_cmd_tag;

  rematch012_in_cmd_accm_inst_kernel_cmd_valid          <= Kernel_inst_rematch012_in_cmd_valid;
  Kernel_inst_rematch012_in_cmd_ready                   <= rematch012_in_cmd_accm_inst_kernel_cmd_ready;
  rematch012_in_cmd_accm_inst_kernel_cmd_firstIdx       <= Kernel_inst_rematch012_in_cmd_firstIdx;
  rematch012_in_cmd_accm_inst_kernel_cmd_lastIdx        <= Kernel_inst_rematch012_in_cmd_lastIdx;
  rematch012_in_cmd_accm_inst_kernel_cmd_tag            <= Kernel_inst_rematch012_in_cmd_tag;

  rematch013_in_cmd_accm_inst_kernel_cmd_valid          <= Kernel_inst_rematch013_in_cmd_valid;
  Kernel_inst_rematch013_in_cmd_ready                   <= rematch013_in_cmd_accm_inst_kernel_cmd_ready;
  rematch013_in_cmd_accm_inst_kernel_cmd_firstIdx       <= Kernel_inst_rematch013_in_cmd_firstIdx;
  rematch013_in_cmd_accm_inst_kernel_cmd_lastIdx        <= Kernel_inst_rematch013_in_cmd_lastIdx;
  rematch013_in_cmd_accm_inst_kernel_cmd_tag            <= Kernel_inst_rematch013_in_cmd_tag;

  rematch014_in_cmd_accm_inst_kernel_cmd_valid          <= Kernel_inst_rematch014_in_cmd_valid;
  Kernel_inst_rematch014_in_cmd_ready                   <= rematch014_in_cmd_accm_inst_kernel_cmd_ready;
  rematch014_in_cmd_accm_inst_kernel_cmd_firstIdx       <= Kernel_inst_rematch014_in_cmd_firstIdx;
  rematch014_in_cmd_accm_inst_kernel_cmd_lastIdx        <= Kernel_inst_rematch014_in_cmd_lastIdx;
  rematch014_in_cmd_accm_inst_kernel_cmd_tag            <= Kernel_inst_rematch014_in_cmd_tag;

  rematch015_in_cmd_accm_inst_kernel_cmd_valid          <= Kernel_inst_rematch015_in_cmd_valid;
  Kernel_inst_rematch015_in_cmd_ready                   <= rematch015_in_cmd_accm_inst_kernel_cmd_ready;
  rematch015_in_cmd_accm_inst_kernel_cmd_firstIdx       <= Kernel_inst_rematch015_in_cmd_firstIdx;
  rematch015_in_cmd_accm_inst_kernel_cmd_lastIdx        <= Kernel_inst_rematch015_in_cmd_lastIdx;
  rematch015_in_cmd_accm_inst_kernel_cmd_tag            <= Kernel_inst_rematch015_in_cmd_tag;

  rematch000_taxi_out_cmd_accm_inst_kernel_cmd_valid    <= Kernel_inst_rematch000_taxi_out_cmd_valid;
  Kernel_inst_rematch000_taxi_out_cmd_ready             <= rematch000_taxi_out_cmd_accm_inst_kernel_cmd_ready;
  rematch000_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx <= Kernel_inst_rematch000_taxi_out_cmd_firstIdx;
  rematch000_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx  <= Kernel_inst_rematch000_taxi_out_cmd_lastIdx;
  rematch000_taxi_out_cmd_accm_inst_kernel_cmd_tag      <= Kernel_inst_rematch000_taxi_out_cmd_tag;

  rematch001_taxi_out_cmd_accm_inst_kernel_cmd_valid    <= Kernel_inst_rematch001_taxi_out_cmd_valid;
  Kernel_inst_rematch001_taxi_out_cmd_ready             <= rematch001_taxi_out_cmd_accm_inst_kernel_cmd_ready;
  rematch001_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx <= Kernel_inst_rematch001_taxi_out_cmd_firstIdx;
  rematch001_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx  <= Kernel_inst_rematch001_taxi_out_cmd_lastIdx;
  rematch001_taxi_out_cmd_accm_inst_kernel_cmd_tag      <= Kernel_inst_rematch001_taxi_out_cmd_tag;

  rematch002_taxi_out_cmd_accm_inst_kernel_cmd_valid    <= Kernel_inst_rematch002_taxi_out_cmd_valid;
  Kernel_inst_rematch002_taxi_out_cmd_ready             <= rematch002_taxi_out_cmd_accm_inst_kernel_cmd_ready;
  rematch002_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx <= Kernel_inst_rematch002_taxi_out_cmd_firstIdx;
  rematch002_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx  <= Kernel_inst_rematch002_taxi_out_cmd_lastIdx;
  rematch002_taxi_out_cmd_accm_inst_kernel_cmd_tag      <= Kernel_inst_rematch002_taxi_out_cmd_tag;

  rematch003_taxi_out_cmd_accm_inst_kernel_cmd_valid    <= Kernel_inst_rematch003_taxi_out_cmd_valid;
  Kernel_inst_rematch003_taxi_out_cmd_ready             <= rematch003_taxi_out_cmd_accm_inst_kernel_cmd_ready;
  rematch003_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx <= Kernel_inst_rematch003_taxi_out_cmd_firstIdx;
  rematch003_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx  <= Kernel_inst_rematch003_taxi_out_cmd_lastIdx;
  rematch003_taxi_out_cmd_accm_inst_kernel_cmd_tag      <= Kernel_inst_rematch003_taxi_out_cmd_tag;

  rematch004_taxi_out_cmd_accm_inst_kernel_cmd_valid    <= Kernel_inst_rematch004_taxi_out_cmd_valid;
  Kernel_inst_rematch004_taxi_out_cmd_ready             <= rematch004_taxi_out_cmd_accm_inst_kernel_cmd_ready;
  rematch004_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx <= Kernel_inst_rematch004_taxi_out_cmd_firstIdx;
  rematch004_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx  <= Kernel_inst_rematch004_taxi_out_cmd_lastIdx;
  rematch004_taxi_out_cmd_accm_inst_kernel_cmd_tag      <= Kernel_inst_rematch004_taxi_out_cmd_tag;

  rematch005_taxi_out_cmd_accm_inst_kernel_cmd_valid    <= Kernel_inst_rematch005_taxi_out_cmd_valid;
  Kernel_inst_rematch005_taxi_out_cmd_ready             <= rematch005_taxi_out_cmd_accm_inst_kernel_cmd_ready;
  rematch005_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx <= Kernel_inst_rematch005_taxi_out_cmd_firstIdx;
  rematch005_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx  <= Kernel_inst_rematch005_taxi_out_cmd_lastIdx;
  rematch005_taxi_out_cmd_accm_inst_kernel_cmd_tag      <= Kernel_inst_rematch005_taxi_out_cmd_tag;

  rematch006_taxi_out_cmd_accm_inst_kernel_cmd_valid    <= Kernel_inst_rematch006_taxi_out_cmd_valid;
  Kernel_inst_rematch006_taxi_out_cmd_ready             <= rematch006_taxi_out_cmd_accm_inst_kernel_cmd_ready;
  rematch006_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx <= Kernel_inst_rematch006_taxi_out_cmd_firstIdx;
  rematch006_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx  <= Kernel_inst_rematch006_taxi_out_cmd_lastIdx;
  rematch006_taxi_out_cmd_accm_inst_kernel_cmd_tag      <= Kernel_inst_rematch006_taxi_out_cmd_tag;

  rematch007_taxi_out_cmd_accm_inst_kernel_cmd_valid    <= Kernel_inst_rematch007_taxi_out_cmd_valid;
  Kernel_inst_rematch007_taxi_out_cmd_ready             <= rematch007_taxi_out_cmd_accm_inst_kernel_cmd_ready;
  rematch007_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx <= Kernel_inst_rematch007_taxi_out_cmd_firstIdx;
  rematch007_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx  <= Kernel_inst_rematch007_taxi_out_cmd_lastIdx;
  rematch007_taxi_out_cmd_accm_inst_kernel_cmd_tag      <= Kernel_inst_rematch007_taxi_out_cmd_tag;

  rematch008_taxi_out_cmd_accm_inst_kernel_cmd_valid    <= Kernel_inst_rematch008_taxi_out_cmd_valid;
  Kernel_inst_rematch008_taxi_out_cmd_ready             <= rematch008_taxi_out_cmd_accm_inst_kernel_cmd_ready;
  rematch008_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx <= Kernel_inst_rematch008_taxi_out_cmd_firstIdx;
  rematch008_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx  <= Kernel_inst_rematch008_taxi_out_cmd_lastIdx;
  rematch008_taxi_out_cmd_accm_inst_kernel_cmd_tag      <= Kernel_inst_rematch008_taxi_out_cmd_tag;

  rematch009_taxi_out_cmd_accm_inst_kernel_cmd_valid    <= Kernel_inst_rematch009_taxi_out_cmd_valid;
  Kernel_inst_rematch009_taxi_out_cmd_ready             <= rematch009_taxi_out_cmd_accm_inst_kernel_cmd_ready;
  rematch009_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx <= Kernel_inst_rematch009_taxi_out_cmd_firstIdx;
  rematch009_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx  <= Kernel_inst_rematch009_taxi_out_cmd_lastIdx;
  rematch009_taxi_out_cmd_accm_inst_kernel_cmd_tag      <= Kernel_inst_rematch009_taxi_out_cmd_tag;

  rematch010_taxi_out_cmd_accm_inst_kernel_cmd_valid    <= Kernel_inst_rematch010_taxi_out_cmd_valid;
  Kernel_inst_rematch010_taxi_out_cmd_ready             <= rematch010_taxi_out_cmd_accm_inst_kernel_cmd_ready;
  rematch010_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx <= Kernel_inst_rematch010_taxi_out_cmd_firstIdx;
  rematch010_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx  <= Kernel_inst_rematch010_taxi_out_cmd_lastIdx;
  rematch010_taxi_out_cmd_accm_inst_kernel_cmd_tag      <= Kernel_inst_rematch010_taxi_out_cmd_tag;

  rematch011_taxi_out_cmd_accm_inst_kernel_cmd_valid    <= Kernel_inst_rematch011_taxi_out_cmd_valid;
  Kernel_inst_rematch011_taxi_out_cmd_ready             <= rematch011_taxi_out_cmd_accm_inst_kernel_cmd_ready;
  rematch011_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx <= Kernel_inst_rematch011_taxi_out_cmd_firstIdx;
  rematch011_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx  <= Kernel_inst_rematch011_taxi_out_cmd_lastIdx;
  rematch011_taxi_out_cmd_accm_inst_kernel_cmd_tag      <= Kernel_inst_rematch011_taxi_out_cmd_tag;

  rematch012_taxi_out_cmd_accm_inst_kernel_cmd_valid    <= Kernel_inst_rematch012_taxi_out_cmd_valid;
  Kernel_inst_rematch012_taxi_out_cmd_ready             <= rematch012_taxi_out_cmd_accm_inst_kernel_cmd_ready;
  rematch012_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx <= Kernel_inst_rematch012_taxi_out_cmd_firstIdx;
  rematch012_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx  <= Kernel_inst_rematch012_taxi_out_cmd_lastIdx;
  rematch012_taxi_out_cmd_accm_inst_kernel_cmd_tag      <= Kernel_inst_rematch012_taxi_out_cmd_tag;

  rematch013_taxi_out_cmd_accm_inst_kernel_cmd_valid    <= Kernel_inst_rematch013_taxi_out_cmd_valid;
  Kernel_inst_rematch013_taxi_out_cmd_ready             <= rematch013_taxi_out_cmd_accm_inst_kernel_cmd_ready;
  rematch013_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx <= Kernel_inst_rematch013_taxi_out_cmd_firstIdx;
  rematch013_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx  <= Kernel_inst_rematch013_taxi_out_cmd_lastIdx;
  rematch013_taxi_out_cmd_accm_inst_kernel_cmd_tag      <= Kernel_inst_rematch013_taxi_out_cmd_tag;

  rematch014_taxi_out_cmd_accm_inst_kernel_cmd_valid    <= Kernel_inst_rematch014_taxi_out_cmd_valid;
  Kernel_inst_rematch014_taxi_out_cmd_ready             <= rematch014_taxi_out_cmd_accm_inst_kernel_cmd_ready;
  rematch014_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx <= Kernel_inst_rematch014_taxi_out_cmd_firstIdx;
  rematch014_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx  <= Kernel_inst_rematch014_taxi_out_cmd_lastIdx;
  rematch014_taxi_out_cmd_accm_inst_kernel_cmd_tag      <= Kernel_inst_rematch014_taxi_out_cmd_tag;

  rematch015_taxi_out_cmd_accm_inst_kernel_cmd_valid    <= Kernel_inst_rematch015_taxi_out_cmd_valid;
  Kernel_inst_rematch015_taxi_out_cmd_ready             <= rematch015_taxi_out_cmd_accm_inst_kernel_cmd_ready;
  rematch015_taxi_out_cmd_accm_inst_kernel_cmd_firstIdx <= Kernel_inst_rematch015_taxi_out_cmd_firstIdx;
  rematch015_taxi_out_cmd_accm_inst_kernel_cmd_lastIdx  <= Kernel_inst_rematch015_taxi_out_cmd_lastIdx;
  rematch015_taxi_out_cmd_accm_inst_kernel_cmd_tag      <= Kernel_inst_rematch015_taxi_out_cmd_tag;

  rematch000_in_cmd_accm_inst_ctrl(63 downto 0)       <= mmio_inst_f_rematch000_in_offsets_data;
  rematch000_in_cmd_accm_inst_ctrl(127 downto 64)     <= mmio_inst_f_rematch000_in_values_data;

  rematch001_in_cmd_accm_inst_ctrl(63 downto 0)       <= mmio_inst_f_rematch001_in_offsets_data;
  rematch001_in_cmd_accm_inst_ctrl(127 downto 64)     <= mmio_inst_f_rematch001_in_values_data;

  rematch002_in_cmd_accm_inst_ctrl(63 downto 0)       <= mmio_inst_f_rematch002_in_offsets_data;
  rematch002_in_cmd_accm_inst_ctrl(127 downto 64)     <= mmio_inst_f_rematch002_in_values_data;

  rematch003_in_cmd_accm_inst_ctrl(63 downto 0)       <= mmio_inst_f_rematch003_in_offsets_data;
  rematch003_in_cmd_accm_inst_ctrl(127 downto 64)     <= mmio_inst_f_rematch003_in_values_data;

  rematch004_in_cmd_accm_inst_ctrl(63 downto 0)       <= mmio_inst_f_rematch004_in_offsets_data;
  rematch004_in_cmd_accm_inst_ctrl(127 downto 64)     <= mmio_inst_f_rematch004_in_values_data;

  rematch005_in_cmd_accm_inst_ctrl(63 downto 0)       <= mmio_inst_f_rematch005_in_offsets_data;
  rematch005_in_cmd_accm_inst_ctrl(127 downto 64)     <= mmio_inst_f_rematch005_in_values_data;

  rematch006_in_cmd_accm_inst_ctrl(63 downto 0)       <= mmio_inst_f_rematch006_in_offsets_data;
  rematch006_in_cmd_accm_inst_ctrl(127 downto 64)     <= mmio_inst_f_rematch006_in_values_data;

  rematch007_in_cmd_accm_inst_ctrl(63 downto 0)       <= mmio_inst_f_rematch007_in_offsets_data;
  rematch007_in_cmd_accm_inst_ctrl(127 downto 64)     <= mmio_inst_f_rematch007_in_values_data;

  rematch008_in_cmd_accm_inst_ctrl(63 downto 0)       <= mmio_inst_f_rematch008_in_offsets_data;
  rematch008_in_cmd_accm_inst_ctrl(127 downto 64)     <= mmio_inst_f_rematch008_in_values_data;

  rematch009_in_cmd_accm_inst_ctrl(63 downto 0)       <= mmio_inst_f_rematch009_in_offsets_data;
  rematch009_in_cmd_accm_inst_ctrl(127 downto 64)     <= mmio_inst_f_rematch009_in_values_data;

  rematch010_in_cmd_accm_inst_ctrl(63 downto 0)       <= mmio_inst_f_rematch010_in_offsets_data;
  rematch010_in_cmd_accm_inst_ctrl(127 downto 64)     <= mmio_inst_f_rematch010_in_values_data;

  rematch011_in_cmd_accm_inst_ctrl(63 downto 0)       <= mmio_inst_f_rematch011_in_offsets_data;
  rematch011_in_cmd_accm_inst_ctrl(127 downto 64)     <= mmio_inst_f_rematch011_in_values_data;

  rematch012_in_cmd_accm_inst_ctrl(63 downto 0)       <= mmio_inst_f_rematch012_in_offsets_data;
  rematch012_in_cmd_accm_inst_ctrl(127 downto 64)     <= mmio_inst_f_rematch012_in_values_data;

  rematch013_in_cmd_accm_inst_ctrl(63 downto 0)       <= mmio_inst_f_rematch013_in_offsets_data;
  rematch013_in_cmd_accm_inst_ctrl(127 downto 64)     <= mmio_inst_f_rematch013_in_values_data;

  rematch014_in_cmd_accm_inst_ctrl(63 downto 0)       <= mmio_inst_f_rematch014_in_offsets_data;
  rematch014_in_cmd_accm_inst_ctrl(127 downto 64)     <= mmio_inst_f_rematch014_in_values_data;

  rematch015_in_cmd_accm_inst_ctrl(63 downto 0)       <= mmio_inst_f_rematch015_in_offsets_data;
  rematch015_in_cmd_accm_inst_ctrl(127 downto 64)     <= mmio_inst_f_rematch015_in_values_data;

  rematch000_taxi_out_cmd_accm_inst_ctrl(63 downto 0) <= mmio_inst_f_rematch000_taxi_out_values_data;
  rematch001_taxi_out_cmd_accm_inst_ctrl(63 downto 0) <= mmio_inst_f_rematch001_taxi_out_values_data;
  rematch002_taxi_out_cmd_accm_inst_ctrl(63 downto 0) <= mmio_inst_f_rematch002_taxi_out_values_data;
  rematch003_taxi_out_cmd_accm_inst_ctrl(63 downto 0) <= mmio_inst_f_rematch003_taxi_out_values_data;
  rematch004_taxi_out_cmd_accm_inst_ctrl(63 downto 0) <= mmio_inst_f_rematch004_taxi_out_values_data;
  rematch005_taxi_out_cmd_accm_inst_ctrl(63 downto 0) <= mmio_inst_f_rematch005_taxi_out_values_data;
  rematch006_taxi_out_cmd_accm_inst_ctrl(63 downto 0) <= mmio_inst_f_rematch006_taxi_out_values_data;
  rematch007_taxi_out_cmd_accm_inst_ctrl(63 downto 0) <= mmio_inst_f_rematch007_taxi_out_values_data;
  rematch008_taxi_out_cmd_accm_inst_ctrl(63 downto 0) <= mmio_inst_f_rematch008_taxi_out_values_data;
  rematch009_taxi_out_cmd_accm_inst_ctrl(63 downto 0) <= mmio_inst_f_rematch009_taxi_out_values_data;
  rematch010_taxi_out_cmd_accm_inst_ctrl(63 downto 0) <= mmio_inst_f_rematch010_taxi_out_values_data;
  rematch011_taxi_out_cmd_accm_inst_ctrl(63 downto 0) <= mmio_inst_f_rematch011_taxi_out_values_data;
  rematch012_taxi_out_cmd_accm_inst_ctrl(63 downto 0) <= mmio_inst_f_rematch012_taxi_out_values_data;
  rematch013_taxi_out_cmd_accm_inst_ctrl(63 downto 0) <= mmio_inst_f_rematch013_taxi_out_values_data;
  rematch014_taxi_out_cmd_accm_inst_ctrl(63 downto 0) <= mmio_inst_f_rematch014_taxi_out_values_data;
  rematch015_taxi_out_cmd_accm_inst_ctrl(63 downto 0) <= mmio_inst_f_rematch015_taxi_out_values_data;

end architecture;
