-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.Interconnect_pkg.all;

entity Kernel_Mantle is
  generic (
    INDEX_WIDTH        : integer := 32;
    TAG_WIDTH          : integer := 1;
    BUS_ADDR_WIDTH     : integer := 64;
    BUS_DATA_WIDTH     : integer := 512;
    BUS_LEN_WIDTH      : integer := 8;
    BUS_BURST_STEP_LEN : integer := 1;
    BUS_BURST_MAX_LEN  : integer := 16
  );
  port (
    bcd_clk           : in  std_logic;
    bcd_reset         : in  std_logic;
    kcd_clk           : in  std_logic;
    kcd_reset         : in  std_logic;
    mmio_awvalid      : in  std_logic;
    mmio_awready      : out std_logic;
    mmio_awaddr       : in  std_logic_vector(31 downto 0);
    mmio_wvalid       : in  std_logic;
    mmio_wready       : out std_logic;
    mmio_wdata        : in  std_logic_vector(31 downto 0);
    mmio_wstrb        : in  std_logic_vector(3 downto 0);
    mmio_bvalid       : out std_logic;
    mmio_bready       : in  std_logic;
    mmio_bresp        : out std_logic_vector(1 downto 0);
    mmio_arvalid      : in  std_logic;
    mmio_arready      : out std_logic;
    mmio_araddr       : in  std_logic_vector(31 downto 0);
    mmio_rvalid       : out std_logic;
    mmio_rready       : in  std_logic;
    mmio_rdata        : out std_logic_vector(31 downto 0);
    mmio_rresp        : out std_logic_vector(1 downto 0);
    rd_mst_rreq_valid : out std_logic;
    rd_mst_rreq_ready : in  std_logic;
    rd_mst_rreq_addr  : out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    rd_mst_rreq_len   : out std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
    rd_mst_rdat_valid : in  std_logic;
    rd_mst_rdat_ready : out std_logic;
    rd_mst_rdat_data  : in  std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
    rd_mst_rdat_last  : in  std_logic
  );
end entity;

architecture Implementation of Kernel_Mantle is
  component Kernel_Nucleus is
    generic (
      INDEX_WIDTH                  : integer := 32;
      TAG_WIDTH                    : integer := 1;
      REMATCH000_IN_BUS_ADDR_WIDTH : integer := 64;
      REMATCH001_IN_BUS_ADDR_WIDTH : integer := 64;
      REMATCH002_IN_BUS_ADDR_WIDTH : integer := 64;
      REMATCH003_IN_BUS_ADDR_WIDTH : integer := 64;
      REMATCH004_IN_BUS_ADDR_WIDTH : integer := 64;
      REMATCH005_IN_BUS_ADDR_WIDTH : integer := 64;
      REMATCH006_IN_BUS_ADDR_WIDTH : integer := 64;
      REMATCH007_IN_BUS_ADDR_WIDTH : integer := 64;
      REMATCH008_IN_BUS_ADDR_WIDTH : integer := 64;
      REMATCH009_IN_BUS_ADDR_WIDTH : integer := 64;
      REMATCH010_IN_BUS_ADDR_WIDTH : integer := 64;
      REMATCH011_IN_BUS_ADDR_WIDTH : integer := 64;
      REMATCH012_IN_BUS_ADDR_WIDTH : integer := 64;
      REMATCH013_IN_BUS_ADDR_WIDTH : integer := 64;
      REMATCH014_IN_BUS_ADDR_WIDTH : integer := 64;
      REMATCH015_IN_BUS_ADDR_WIDTH : integer := 64
    );
    port (
      kcd_clk                    : in  std_logic;
      kcd_reset                  : in  std_logic;
      mmio_awvalid               : in  std_logic;
      mmio_awready               : out std_logic;
      mmio_awaddr                : in  std_logic_vector(31 downto 0);
      mmio_wvalid                : in  std_logic;
      mmio_wready                : out std_logic;
      mmio_wdata                 : in  std_logic_vector(31 downto 0);
      mmio_wstrb                 : in  std_logic_vector(3 downto 0);
      mmio_bvalid                : out std_logic;
      mmio_bready                : in  std_logic;
      mmio_bresp                 : out std_logic_vector(1 downto 0);
      mmio_arvalid               : in  std_logic;
      mmio_arready               : out std_logic;
      mmio_araddr                : in  std_logic_vector(31 downto 0);
      mmio_rvalid                : out std_logic;
      mmio_rready                : in  std_logic;
      mmio_rdata                 : out std_logic_vector(31 downto 0);
      mmio_rresp                 : out std_logic_vector(1 downto 0);
      rematch000_in_valid        : in  std_logic;
      rematch000_in_ready        : out std_logic;
      rematch000_in_dvalid       : in  std_logic;
      rematch000_in_last         : in  std_logic;
      rematch000_in_length       : in  std_logic_vector(31 downto 0);
      rematch000_in_count        : in  std_logic_vector(0 downto 0);
      rematch000_in_chars_valid  : in  std_logic;
      rematch000_in_chars_ready  : out std_logic;
      rematch000_in_chars_dvalid : in  std_logic;
      rematch000_in_chars_last   : in  std_logic;
      rematch000_in_chars        : in  std_logic_vector(31 downto 0);
      rematch000_in_chars_count  : in  std_logic_vector(2 downto 0);
      rematch000_in_unl_valid    : in  std_logic;
      rematch000_in_unl_ready    : out std_logic;
      rematch000_in_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch000_in_cmd_valid    : out std_logic;
      rematch000_in_cmd_ready    : in  std_logic;
      rematch000_in_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch000_in_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch000_in_cmd_ctrl     : out std_logic_vector(REMATCH000_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch000_in_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch001_in_valid        : in  std_logic;
      rematch001_in_ready        : out std_logic;
      rematch001_in_dvalid       : in  std_logic;
      rematch001_in_last         : in  std_logic;
      rematch001_in_length       : in  std_logic_vector(31 downto 0);
      rematch001_in_count        : in  std_logic_vector(0 downto 0);
      rematch001_in_chars_valid  : in  std_logic;
      rematch001_in_chars_ready  : out std_logic;
      rematch001_in_chars_dvalid : in  std_logic;
      rematch001_in_chars_last   : in  std_logic;
      rematch001_in_chars        : in  std_logic_vector(31 downto 0);
      rematch001_in_chars_count  : in  std_logic_vector(2 downto 0);
      rematch001_in_unl_valid    : in  std_logic;
      rematch001_in_unl_ready    : out std_logic;
      rematch001_in_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch001_in_cmd_valid    : out std_logic;
      rematch001_in_cmd_ready    : in  std_logic;
      rematch001_in_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch001_in_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch001_in_cmd_ctrl     : out std_logic_vector(REMATCH001_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch001_in_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch002_in_valid        : in  std_logic;
      rematch002_in_ready        : out std_logic;
      rematch002_in_dvalid       : in  std_logic;
      rematch002_in_last         : in  std_logic;
      rematch002_in_length       : in  std_logic_vector(31 downto 0);
      rematch002_in_count        : in  std_logic_vector(0 downto 0);
      rematch002_in_chars_valid  : in  std_logic;
      rematch002_in_chars_ready  : out std_logic;
      rematch002_in_chars_dvalid : in  std_logic;
      rematch002_in_chars_last   : in  std_logic;
      rematch002_in_chars        : in  std_logic_vector(31 downto 0);
      rematch002_in_chars_count  : in  std_logic_vector(2 downto 0);
      rematch002_in_unl_valid    : in  std_logic;
      rematch002_in_unl_ready    : out std_logic;
      rematch002_in_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch002_in_cmd_valid    : out std_logic;
      rematch002_in_cmd_ready    : in  std_logic;
      rematch002_in_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch002_in_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch002_in_cmd_ctrl     : out std_logic_vector(REMATCH002_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch002_in_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch003_in_valid        : in  std_logic;
      rematch003_in_ready        : out std_logic;
      rematch003_in_dvalid       : in  std_logic;
      rematch003_in_last         : in  std_logic;
      rematch003_in_length       : in  std_logic_vector(31 downto 0);
      rematch003_in_count        : in  std_logic_vector(0 downto 0);
      rematch003_in_chars_valid  : in  std_logic;
      rematch003_in_chars_ready  : out std_logic;
      rematch003_in_chars_dvalid : in  std_logic;
      rematch003_in_chars_last   : in  std_logic;
      rematch003_in_chars        : in  std_logic_vector(31 downto 0);
      rematch003_in_chars_count  : in  std_logic_vector(2 downto 0);
      rematch003_in_unl_valid    : in  std_logic;
      rematch003_in_unl_ready    : out std_logic;
      rematch003_in_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch003_in_cmd_valid    : out std_logic;
      rematch003_in_cmd_ready    : in  std_logic;
      rematch003_in_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch003_in_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch003_in_cmd_ctrl     : out std_logic_vector(REMATCH003_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch003_in_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch004_in_valid        : in  std_logic;
      rematch004_in_ready        : out std_logic;
      rematch004_in_dvalid       : in  std_logic;
      rematch004_in_last         : in  std_logic;
      rematch004_in_length       : in  std_logic_vector(31 downto 0);
      rematch004_in_count        : in  std_logic_vector(0 downto 0);
      rematch004_in_chars_valid  : in  std_logic;
      rematch004_in_chars_ready  : out std_logic;
      rematch004_in_chars_dvalid : in  std_logic;
      rematch004_in_chars_last   : in  std_logic;
      rematch004_in_chars        : in  std_logic_vector(31 downto 0);
      rematch004_in_chars_count  : in  std_logic_vector(2 downto 0);
      rematch004_in_unl_valid    : in  std_logic;
      rematch004_in_unl_ready    : out std_logic;
      rematch004_in_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch004_in_cmd_valid    : out std_logic;
      rematch004_in_cmd_ready    : in  std_logic;
      rematch004_in_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch004_in_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch004_in_cmd_ctrl     : out std_logic_vector(REMATCH004_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch004_in_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch005_in_valid        : in  std_logic;
      rematch005_in_ready        : out std_logic;
      rematch005_in_dvalid       : in  std_logic;
      rematch005_in_last         : in  std_logic;
      rematch005_in_length       : in  std_logic_vector(31 downto 0);
      rematch005_in_count        : in  std_logic_vector(0 downto 0);
      rematch005_in_chars_valid  : in  std_logic;
      rematch005_in_chars_ready  : out std_logic;
      rematch005_in_chars_dvalid : in  std_logic;
      rematch005_in_chars_last   : in  std_logic;
      rematch005_in_chars        : in  std_logic_vector(31 downto 0);
      rematch005_in_chars_count  : in  std_logic_vector(2 downto 0);
      rematch005_in_unl_valid    : in  std_logic;
      rematch005_in_unl_ready    : out std_logic;
      rematch005_in_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch005_in_cmd_valid    : out std_logic;
      rematch005_in_cmd_ready    : in  std_logic;
      rematch005_in_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch005_in_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch005_in_cmd_ctrl     : out std_logic_vector(REMATCH005_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch005_in_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch006_in_valid        : in  std_logic;
      rematch006_in_ready        : out std_logic;
      rematch006_in_dvalid       : in  std_logic;
      rematch006_in_last         : in  std_logic;
      rematch006_in_length       : in  std_logic_vector(31 downto 0);
      rematch006_in_count        : in  std_logic_vector(0 downto 0);
      rematch006_in_chars_valid  : in  std_logic;
      rematch006_in_chars_ready  : out std_logic;
      rematch006_in_chars_dvalid : in  std_logic;
      rematch006_in_chars_last   : in  std_logic;
      rematch006_in_chars        : in  std_logic_vector(31 downto 0);
      rematch006_in_chars_count  : in  std_logic_vector(2 downto 0);
      rematch006_in_unl_valid    : in  std_logic;
      rematch006_in_unl_ready    : out std_logic;
      rematch006_in_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch006_in_cmd_valid    : out std_logic;
      rematch006_in_cmd_ready    : in  std_logic;
      rematch006_in_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch006_in_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch006_in_cmd_ctrl     : out std_logic_vector(REMATCH006_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch006_in_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch007_in_valid        : in  std_logic;
      rematch007_in_ready        : out std_logic;
      rematch007_in_dvalid       : in  std_logic;
      rematch007_in_last         : in  std_logic;
      rematch007_in_length       : in  std_logic_vector(31 downto 0);
      rematch007_in_count        : in  std_logic_vector(0 downto 0);
      rematch007_in_chars_valid  : in  std_logic;
      rematch007_in_chars_ready  : out std_logic;
      rematch007_in_chars_dvalid : in  std_logic;
      rematch007_in_chars_last   : in  std_logic;
      rematch007_in_chars        : in  std_logic_vector(31 downto 0);
      rematch007_in_chars_count  : in  std_logic_vector(2 downto 0);
      rematch007_in_unl_valid    : in  std_logic;
      rematch007_in_unl_ready    : out std_logic;
      rematch007_in_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch007_in_cmd_valid    : out std_logic;
      rematch007_in_cmd_ready    : in  std_logic;
      rematch007_in_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch007_in_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch007_in_cmd_ctrl     : out std_logic_vector(REMATCH007_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch007_in_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch008_in_valid        : in  std_logic;
      rematch008_in_ready        : out std_logic;
      rematch008_in_dvalid       : in  std_logic;
      rematch008_in_last         : in  std_logic;
      rematch008_in_length       : in  std_logic_vector(31 downto 0);
      rematch008_in_count        : in  std_logic_vector(0 downto 0);
      rematch008_in_chars_valid  : in  std_logic;
      rematch008_in_chars_ready  : out std_logic;
      rematch008_in_chars_dvalid : in  std_logic;
      rematch008_in_chars_last   : in  std_logic;
      rematch008_in_chars        : in  std_logic_vector(31 downto 0);
      rematch008_in_chars_count  : in  std_logic_vector(2 downto 0);
      rematch008_in_unl_valid    : in  std_logic;
      rematch008_in_unl_ready    : out std_logic;
      rematch008_in_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch008_in_cmd_valid    : out std_logic;
      rematch008_in_cmd_ready    : in  std_logic;
      rematch008_in_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch008_in_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch008_in_cmd_ctrl     : out std_logic_vector(REMATCH008_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch008_in_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch009_in_valid        : in  std_logic;
      rematch009_in_ready        : out std_logic;
      rematch009_in_dvalid       : in  std_logic;
      rematch009_in_last         : in  std_logic;
      rematch009_in_length       : in  std_logic_vector(31 downto 0);
      rematch009_in_count        : in  std_logic_vector(0 downto 0);
      rematch009_in_chars_valid  : in  std_logic;
      rematch009_in_chars_ready  : out std_logic;
      rematch009_in_chars_dvalid : in  std_logic;
      rematch009_in_chars_last   : in  std_logic;
      rematch009_in_chars        : in  std_logic_vector(31 downto 0);
      rematch009_in_chars_count  : in  std_logic_vector(2 downto 0);
      rematch009_in_unl_valid    : in  std_logic;
      rematch009_in_unl_ready    : out std_logic;
      rematch009_in_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch009_in_cmd_valid    : out std_logic;
      rematch009_in_cmd_ready    : in  std_logic;
      rematch009_in_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch009_in_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch009_in_cmd_ctrl     : out std_logic_vector(REMATCH009_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch009_in_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch010_in_valid        : in  std_logic;
      rematch010_in_ready        : out std_logic;
      rematch010_in_dvalid       : in  std_logic;
      rematch010_in_last         : in  std_logic;
      rematch010_in_length       : in  std_logic_vector(31 downto 0);
      rematch010_in_count        : in  std_logic_vector(0 downto 0);
      rematch010_in_chars_valid  : in  std_logic;
      rematch010_in_chars_ready  : out std_logic;
      rematch010_in_chars_dvalid : in  std_logic;
      rematch010_in_chars_last   : in  std_logic;
      rematch010_in_chars        : in  std_logic_vector(31 downto 0);
      rematch010_in_chars_count  : in  std_logic_vector(2 downto 0);
      rematch010_in_unl_valid    : in  std_logic;
      rematch010_in_unl_ready    : out std_logic;
      rematch010_in_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch010_in_cmd_valid    : out std_logic;
      rematch010_in_cmd_ready    : in  std_logic;
      rematch010_in_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch010_in_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch010_in_cmd_ctrl     : out std_logic_vector(REMATCH010_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch010_in_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch011_in_valid        : in  std_logic;
      rematch011_in_ready        : out std_logic;
      rematch011_in_dvalid       : in  std_logic;
      rematch011_in_last         : in  std_logic;
      rematch011_in_length       : in  std_logic_vector(31 downto 0);
      rematch011_in_count        : in  std_logic_vector(0 downto 0);
      rematch011_in_chars_valid  : in  std_logic;
      rematch011_in_chars_ready  : out std_logic;
      rematch011_in_chars_dvalid : in  std_logic;
      rematch011_in_chars_last   : in  std_logic;
      rematch011_in_chars        : in  std_logic_vector(31 downto 0);
      rematch011_in_chars_count  : in  std_logic_vector(2 downto 0);
      rematch011_in_unl_valid    : in  std_logic;
      rematch011_in_unl_ready    : out std_logic;
      rematch011_in_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch011_in_cmd_valid    : out std_logic;
      rematch011_in_cmd_ready    : in  std_logic;
      rematch011_in_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch011_in_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch011_in_cmd_ctrl     : out std_logic_vector(REMATCH011_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch011_in_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch012_in_valid        : in  std_logic;
      rematch012_in_ready        : out std_logic;
      rematch012_in_dvalid       : in  std_logic;
      rematch012_in_last         : in  std_logic;
      rematch012_in_length       : in  std_logic_vector(31 downto 0);
      rematch012_in_count        : in  std_logic_vector(0 downto 0);
      rematch012_in_chars_valid  : in  std_logic;
      rematch012_in_chars_ready  : out std_logic;
      rematch012_in_chars_dvalid : in  std_logic;
      rematch012_in_chars_last   : in  std_logic;
      rematch012_in_chars        : in  std_logic_vector(31 downto 0);
      rematch012_in_chars_count  : in  std_logic_vector(2 downto 0);
      rematch012_in_unl_valid    : in  std_logic;
      rematch012_in_unl_ready    : out std_logic;
      rematch012_in_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch012_in_cmd_valid    : out std_logic;
      rematch012_in_cmd_ready    : in  std_logic;
      rematch012_in_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch012_in_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch012_in_cmd_ctrl     : out std_logic_vector(REMATCH012_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch012_in_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch013_in_valid        : in  std_logic;
      rematch013_in_ready        : out std_logic;
      rematch013_in_dvalid       : in  std_logic;
      rematch013_in_last         : in  std_logic;
      rematch013_in_length       : in  std_logic_vector(31 downto 0);
      rematch013_in_count        : in  std_logic_vector(0 downto 0);
      rematch013_in_chars_valid  : in  std_logic;
      rematch013_in_chars_ready  : out std_logic;
      rematch013_in_chars_dvalid : in  std_logic;
      rematch013_in_chars_last   : in  std_logic;
      rematch013_in_chars        : in  std_logic_vector(31 downto 0);
      rematch013_in_chars_count  : in  std_logic_vector(2 downto 0);
      rematch013_in_unl_valid    : in  std_logic;
      rematch013_in_unl_ready    : out std_logic;
      rematch013_in_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch013_in_cmd_valid    : out std_logic;
      rematch013_in_cmd_ready    : in  std_logic;
      rematch013_in_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch013_in_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch013_in_cmd_ctrl     : out std_logic_vector(REMATCH013_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch013_in_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch014_in_valid        : in  std_logic;
      rematch014_in_ready        : out std_logic;
      rematch014_in_dvalid       : in  std_logic;
      rematch014_in_last         : in  std_logic;
      rematch014_in_length       : in  std_logic_vector(31 downto 0);
      rematch014_in_count        : in  std_logic_vector(0 downto 0);
      rematch014_in_chars_valid  : in  std_logic;
      rematch014_in_chars_ready  : out std_logic;
      rematch014_in_chars_dvalid : in  std_logic;
      rematch014_in_chars_last   : in  std_logic;
      rematch014_in_chars        : in  std_logic_vector(31 downto 0);
      rematch014_in_chars_count  : in  std_logic_vector(2 downto 0);
      rematch014_in_unl_valid    : in  std_logic;
      rematch014_in_unl_ready    : out std_logic;
      rematch014_in_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch014_in_cmd_valid    : out std_logic;
      rematch014_in_cmd_ready    : in  std_logic;
      rematch014_in_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch014_in_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch014_in_cmd_ctrl     : out std_logic_vector(REMATCH014_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch014_in_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch015_in_valid        : in  std_logic;
      rematch015_in_ready        : out std_logic;
      rematch015_in_dvalid       : in  std_logic;
      rematch015_in_last         : in  std_logic;
      rematch015_in_length       : in  std_logic_vector(31 downto 0);
      rematch015_in_count        : in  std_logic_vector(0 downto 0);
      rematch015_in_chars_valid  : in  std_logic;
      rematch015_in_chars_ready  : out std_logic;
      rematch015_in_chars_dvalid : in  std_logic;
      rematch015_in_chars_last   : in  std_logic;
      rematch015_in_chars        : in  std_logic_vector(31 downto 0);
      rematch015_in_chars_count  : in  std_logic_vector(2 downto 0);
      rematch015_in_unl_valid    : in  std_logic;
      rematch015_in_unl_ready    : out std_logic;
      rematch015_in_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch015_in_cmd_valid    : out std_logic;
      rematch015_in_cmd_ready    : in  std_logic;
      rematch015_in_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch015_in_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch015_in_cmd_ctrl     : out std_logic_vector(REMATCH015_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch015_in_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  component Kernel_rematch000 is
    generic (
      INDEX_WIDTH                      : integer := 32;
      TAG_WIDTH                        : integer := 1;
      REMATCH000_IN_BUS_ADDR_WIDTH     : integer := 64;
      REMATCH000_IN_BUS_DATA_WIDTH     : integer := 512;
      REMATCH000_IN_BUS_LEN_WIDTH      : integer := 8;
      REMATCH000_IN_BUS_BURST_STEP_LEN : integer := 1;
      REMATCH000_IN_BUS_BURST_MAX_LEN  : integer := 16
    );
    port (
      bcd_clk                      : in  std_logic;
      bcd_reset                    : in  std_logic;
      kcd_clk                      : in  std_logic;
      kcd_reset                    : in  std_logic;
      rematch000_in_valid          : out std_logic;
      rematch000_in_ready          : in  std_logic;
      rematch000_in_dvalid         : out std_logic;
      rematch000_in_last           : out std_logic;
      rematch000_in_length         : out std_logic_vector(31 downto 0);
      rematch000_in_count          : out std_logic_vector(0 downto 0);
      rematch000_in_chars_valid    : out std_logic;
      rematch000_in_chars_ready    : in  std_logic;
      rematch000_in_chars_dvalid   : out std_logic;
      rematch000_in_chars_last     : out std_logic;
      rematch000_in_chars          : out std_logic_vector(31 downto 0);
      rematch000_in_chars_count    : out std_logic_vector(2 downto 0);
      rematch000_in_bus_rreq_valid : out std_logic;
      rematch000_in_bus_rreq_ready : in  std_logic;
      rematch000_in_bus_rreq_addr  : out std_logic_vector(REMATCH000_IN_BUS_ADDR_WIDTH-1 downto 0);
      rematch000_in_bus_rreq_len   : out std_logic_vector(REMATCH000_IN_BUS_LEN_WIDTH-1 downto 0);
      rematch000_in_bus_rdat_valid : in  std_logic;
      rematch000_in_bus_rdat_ready : out std_logic;
      rematch000_in_bus_rdat_data  : in  std_logic_vector(REMATCH000_IN_BUS_DATA_WIDTH-1 downto 0);
      rematch000_in_bus_rdat_last  : in  std_logic;
      rematch000_in_cmd_valid      : in  std_logic;
      rematch000_in_cmd_ready      : out std_logic;
      rematch000_in_cmd_firstIdx   : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch000_in_cmd_lastIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch000_in_cmd_ctrl       : in  std_logic_vector(REMATCH000_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch000_in_cmd_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch000_in_unl_valid      : out std_logic;
      rematch000_in_unl_ready      : in  std_logic;
      rematch000_in_unl_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  component Kernel_rematch001 is
    generic (
      INDEX_WIDTH                      : integer := 32;
      TAG_WIDTH                        : integer := 1;
      REMATCH001_IN_BUS_ADDR_WIDTH     : integer := 64;
      REMATCH001_IN_BUS_DATA_WIDTH     : integer := 512;
      REMATCH001_IN_BUS_LEN_WIDTH      : integer := 8;
      REMATCH001_IN_BUS_BURST_STEP_LEN : integer := 1;
      REMATCH001_IN_BUS_BURST_MAX_LEN  : integer := 16
    );
    port (
      bcd_clk                      : in  std_logic;
      bcd_reset                    : in  std_logic;
      kcd_clk                      : in  std_logic;
      kcd_reset                    : in  std_logic;
      rematch001_in_valid          : out std_logic;
      rematch001_in_ready          : in  std_logic;
      rematch001_in_dvalid         : out std_logic;
      rematch001_in_last           : out std_logic;
      rematch001_in_length         : out std_logic_vector(31 downto 0);
      rematch001_in_count          : out std_logic_vector(0 downto 0);
      rematch001_in_chars_valid    : out std_logic;
      rematch001_in_chars_ready    : in  std_logic;
      rematch001_in_chars_dvalid   : out std_logic;
      rematch001_in_chars_last     : out std_logic;
      rematch001_in_chars          : out std_logic_vector(31 downto 0);
      rematch001_in_chars_count    : out std_logic_vector(2 downto 0);
      rematch001_in_bus_rreq_valid : out std_logic;
      rematch001_in_bus_rreq_ready : in  std_logic;
      rematch001_in_bus_rreq_addr  : out std_logic_vector(REMATCH001_IN_BUS_ADDR_WIDTH-1 downto 0);
      rematch001_in_bus_rreq_len   : out std_logic_vector(REMATCH001_IN_BUS_LEN_WIDTH-1 downto 0);
      rematch001_in_bus_rdat_valid : in  std_logic;
      rematch001_in_bus_rdat_ready : out std_logic;
      rematch001_in_bus_rdat_data  : in  std_logic_vector(REMATCH001_IN_BUS_DATA_WIDTH-1 downto 0);
      rematch001_in_bus_rdat_last  : in  std_logic;
      rematch001_in_cmd_valid      : in  std_logic;
      rematch001_in_cmd_ready      : out std_logic;
      rematch001_in_cmd_firstIdx   : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch001_in_cmd_lastIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch001_in_cmd_ctrl       : in  std_logic_vector(REMATCH001_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch001_in_cmd_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch001_in_unl_valid      : out std_logic;
      rematch001_in_unl_ready      : in  std_logic;
      rematch001_in_unl_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  component Kernel_rematch002 is
    generic (
      INDEX_WIDTH                      : integer := 32;
      TAG_WIDTH                        : integer := 1;
      REMATCH002_IN_BUS_ADDR_WIDTH     : integer := 64;
      REMATCH002_IN_BUS_DATA_WIDTH     : integer := 512;
      REMATCH002_IN_BUS_LEN_WIDTH      : integer := 8;
      REMATCH002_IN_BUS_BURST_STEP_LEN : integer := 1;
      REMATCH002_IN_BUS_BURST_MAX_LEN  : integer := 16
    );
    port (
      bcd_clk                      : in  std_logic;
      bcd_reset                    : in  std_logic;
      kcd_clk                      : in  std_logic;
      kcd_reset                    : in  std_logic;
      rematch002_in_valid          : out std_logic;
      rematch002_in_ready          : in  std_logic;
      rematch002_in_dvalid         : out std_logic;
      rematch002_in_last           : out std_logic;
      rematch002_in_length         : out std_logic_vector(31 downto 0);
      rematch002_in_count          : out std_logic_vector(0 downto 0);
      rematch002_in_chars_valid    : out std_logic;
      rematch002_in_chars_ready    : in  std_logic;
      rematch002_in_chars_dvalid   : out std_logic;
      rematch002_in_chars_last     : out std_logic;
      rematch002_in_chars          : out std_logic_vector(31 downto 0);
      rematch002_in_chars_count    : out std_logic_vector(2 downto 0);
      rematch002_in_bus_rreq_valid : out std_logic;
      rematch002_in_bus_rreq_ready : in  std_logic;
      rematch002_in_bus_rreq_addr  : out std_logic_vector(REMATCH002_IN_BUS_ADDR_WIDTH-1 downto 0);
      rematch002_in_bus_rreq_len   : out std_logic_vector(REMATCH002_IN_BUS_LEN_WIDTH-1 downto 0);
      rematch002_in_bus_rdat_valid : in  std_logic;
      rematch002_in_bus_rdat_ready : out std_logic;
      rematch002_in_bus_rdat_data  : in  std_logic_vector(REMATCH002_IN_BUS_DATA_WIDTH-1 downto 0);
      rematch002_in_bus_rdat_last  : in  std_logic;
      rematch002_in_cmd_valid      : in  std_logic;
      rematch002_in_cmd_ready      : out std_logic;
      rematch002_in_cmd_firstIdx   : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch002_in_cmd_lastIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch002_in_cmd_ctrl       : in  std_logic_vector(REMATCH002_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch002_in_cmd_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch002_in_unl_valid      : out std_logic;
      rematch002_in_unl_ready      : in  std_logic;
      rematch002_in_unl_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  component Kernel_rematch003 is
    generic (
      INDEX_WIDTH                      : integer := 32;
      TAG_WIDTH                        : integer := 1;
      REMATCH003_IN_BUS_ADDR_WIDTH     : integer := 64;
      REMATCH003_IN_BUS_DATA_WIDTH     : integer := 512;
      REMATCH003_IN_BUS_LEN_WIDTH      : integer := 8;
      REMATCH003_IN_BUS_BURST_STEP_LEN : integer := 1;
      REMATCH003_IN_BUS_BURST_MAX_LEN  : integer := 16
    );
    port (
      bcd_clk                      : in  std_logic;
      bcd_reset                    : in  std_logic;
      kcd_clk                      : in  std_logic;
      kcd_reset                    : in  std_logic;
      rematch003_in_valid          : out std_logic;
      rematch003_in_ready          : in  std_logic;
      rematch003_in_dvalid         : out std_logic;
      rematch003_in_last           : out std_logic;
      rematch003_in_length         : out std_logic_vector(31 downto 0);
      rematch003_in_count          : out std_logic_vector(0 downto 0);
      rematch003_in_chars_valid    : out std_logic;
      rematch003_in_chars_ready    : in  std_logic;
      rematch003_in_chars_dvalid   : out std_logic;
      rematch003_in_chars_last     : out std_logic;
      rematch003_in_chars          : out std_logic_vector(31 downto 0);
      rematch003_in_chars_count    : out std_logic_vector(2 downto 0);
      rematch003_in_bus_rreq_valid : out std_logic;
      rematch003_in_bus_rreq_ready : in  std_logic;
      rematch003_in_bus_rreq_addr  : out std_logic_vector(REMATCH003_IN_BUS_ADDR_WIDTH-1 downto 0);
      rematch003_in_bus_rreq_len   : out std_logic_vector(REMATCH003_IN_BUS_LEN_WIDTH-1 downto 0);
      rematch003_in_bus_rdat_valid : in  std_logic;
      rematch003_in_bus_rdat_ready : out std_logic;
      rematch003_in_bus_rdat_data  : in  std_logic_vector(REMATCH003_IN_BUS_DATA_WIDTH-1 downto 0);
      rematch003_in_bus_rdat_last  : in  std_logic;
      rematch003_in_cmd_valid      : in  std_logic;
      rematch003_in_cmd_ready      : out std_logic;
      rematch003_in_cmd_firstIdx   : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch003_in_cmd_lastIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch003_in_cmd_ctrl       : in  std_logic_vector(REMATCH003_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch003_in_cmd_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch003_in_unl_valid      : out std_logic;
      rematch003_in_unl_ready      : in  std_logic;
      rematch003_in_unl_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  component Kernel_rematch004 is
    generic (
      INDEX_WIDTH                      : integer := 32;
      TAG_WIDTH                        : integer := 1;
      REMATCH004_IN_BUS_ADDR_WIDTH     : integer := 64;
      REMATCH004_IN_BUS_DATA_WIDTH     : integer := 512;
      REMATCH004_IN_BUS_LEN_WIDTH      : integer := 8;
      REMATCH004_IN_BUS_BURST_STEP_LEN : integer := 1;
      REMATCH004_IN_BUS_BURST_MAX_LEN  : integer := 16
    );
    port (
      bcd_clk                      : in  std_logic;
      bcd_reset                    : in  std_logic;
      kcd_clk                      : in  std_logic;
      kcd_reset                    : in  std_logic;
      rematch004_in_valid          : out std_logic;
      rematch004_in_ready          : in  std_logic;
      rematch004_in_dvalid         : out std_logic;
      rematch004_in_last           : out std_logic;
      rematch004_in_length         : out std_logic_vector(31 downto 0);
      rematch004_in_count          : out std_logic_vector(0 downto 0);
      rematch004_in_chars_valid    : out std_logic;
      rematch004_in_chars_ready    : in  std_logic;
      rematch004_in_chars_dvalid   : out std_logic;
      rematch004_in_chars_last     : out std_logic;
      rematch004_in_chars          : out std_logic_vector(31 downto 0);
      rematch004_in_chars_count    : out std_logic_vector(2 downto 0);
      rematch004_in_bus_rreq_valid : out std_logic;
      rematch004_in_bus_rreq_ready : in  std_logic;
      rematch004_in_bus_rreq_addr  : out std_logic_vector(REMATCH004_IN_BUS_ADDR_WIDTH-1 downto 0);
      rematch004_in_bus_rreq_len   : out std_logic_vector(REMATCH004_IN_BUS_LEN_WIDTH-1 downto 0);
      rematch004_in_bus_rdat_valid : in  std_logic;
      rematch004_in_bus_rdat_ready : out std_logic;
      rematch004_in_bus_rdat_data  : in  std_logic_vector(REMATCH004_IN_BUS_DATA_WIDTH-1 downto 0);
      rematch004_in_bus_rdat_last  : in  std_logic;
      rematch004_in_cmd_valid      : in  std_logic;
      rematch004_in_cmd_ready      : out std_logic;
      rematch004_in_cmd_firstIdx   : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch004_in_cmd_lastIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch004_in_cmd_ctrl       : in  std_logic_vector(REMATCH004_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch004_in_cmd_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch004_in_unl_valid      : out std_logic;
      rematch004_in_unl_ready      : in  std_logic;
      rematch004_in_unl_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  component Kernel_rematch005 is
    generic (
      INDEX_WIDTH                      : integer := 32;
      TAG_WIDTH                        : integer := 1;
      REMATCH005_IN_BUS_ADDR_WIDTH     : integer := 64;
      REMATCH005_IN_BUS_DATA_WIDTH     : integer := 512;
      REMATCH005_IN_BUS_LEN_WIDTH      : integer := 8;
      REMATCH005_IN_BUS_BURST_STEP_LEN : integer := 1;
      REMATCH005_IN_BUS_BURST_MAX_LEN  : integer := 16
    );
    port (
      bcd_clk                      : in  std_logic;
      bcd_reset                    : in  std_logic;
      kcd_clk                      : in  std_logic;
      kcd_reset                    : in  std_logic;
      rematch005_in_valid          : out std_logic;
      rematch005_in_ready          : in  std_logic;
      rematch005_in_dvalid         : out std_logic;
      rematch005_in_last           : out std_logic;
      rematch005_in_length         : out std_logic_vector(31 downto 0);
      rematch005_in_count          : out std_logic_vector(0 downto 0);
      rematch005_in_chars_valid    : out std_logic;
      rematch005_in_chars_ready    : in  std_logic;
      rematch005_in_chars_dvalid   : out std_logic;
      rematch005_in_chars_last     : out std_logic;
      rematch005_in_chars          : out std_logic_vector(31 downto 0);
      rematch005_in_chars_count    : out std_logic_vector(2 downto 0);
      rematch005_in_bus_rreq_valid : out std_logic;
      rematch005_in_bus_rreq_ready : in  std_logic;
      rematch005_in_bus_rreq_addr  : out std_logic_vector(REMATCH005_IN_BUS_ADDR_WIDTH-1 downto 0);
      rematch005_in_bus_rreq_len   : out std_logic_vector(REMATCH005_IN_BUS_LEN_WIDTH-1 downto 0);
      rematch005_in_bus_rdat_valid : in  std_logic;
      rematch005_in_bus_rdat_ready : out std_logic;
      rematch005_in_bus_rdat_data  : in  std_logic_vector(REMATCH005_IN_BUS_DATA_WIDTH-1 downto 0);
      rematch005_in_bus_rdat_last  : in  std_logic;
      rematch005_in_cmd_valid      : in  std_logic;
      rematch005_in_cmd_ready      : out std_logic;
      rematch005_in_cmd_firstIdx   : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch005_in_cmd_lastIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch005_in_cmd_ctrl       : in  std_logic_vector(REMATCH005_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch005_in_cmd_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch005_in_unl_valid      : out std_logic;
      rematch005_in_unl_ready      : in  std_logic;
      rematch005_in_unl_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  component Kernel_rematch006 is
    generic (
      INDEX_WIDTH                      : integer := 32;
      TAG_WIDTH                        : integer := 1;
      REMATCH006_IN_BUS_ADDR_WIDTH     : integer := 64;
      REMATCH006_IN_BUS_DATA_WIDTH     : integer := 512;
      REMATCH006_IN_BUS_LEN_WIDTH      : integer := 8;
      REMATCH006_IN_BUS_BURST_STEP_LEN : integer := 1;
      REMATCH006_IN_BUS_BURST_MAX_LEN  : integer := 16
    );
    port (
      bcd_clk                      : in  std_logic;
      bcd_reset                    : in  std_logic;
      kcd_clk                      : in  std_logic;
      kcd_reset                    : in  std_logic;
      rematch006_in_valid          : out std_logic;
      rematch006_in_ready          : in  std_logic;
      rematch006_in_dvalid         : out std_logic;
      rematch006_in_last           : out std_logic;
      rematch006_in_length         : out std_logic_vector(31 downto 0);
      rematch006_in_count          : out std_logic_vector(0 downto 0);
      rematch006_in_chars_valid    : out std_logic;
      rematch006_in_chars_ready    : in  std_logic;
      rematch006_in_chars_dvalid   : out std_logic;
      rematch006_in_chars_last     : out std_logic;
      rematch006_in_chars          : out std_logic_vector(31 downto 0);
      rematch006_in_chars_count    : out std_logic_vector(2 downto 0);
      rematch006_in_bus_rreq_valid : out std_logic;
      rematch006_in_bus_rreq_ready : in  std_logic;
      rematch006_in_bus_rreq_addr  : out std_logic_vector(REMATCH006_IN_BUS_ADDR_WIDTH-1 downto 0);
      rematch006_in_bus_rreq_len   : out std_logic_vector(REMATCH006_IN_BUS_LEN_WIDTH-1 downto 0);
      rematch006_in_bus_rdat_valid : in  std_logic;
      rematch006_in_bus_rdat_ready : out std_logic;
      rematch006_in_bus_rdat_data  : in  std_logic_vector(REMATCH006_IN_BUS_DATA_WIDTH-1 downto 0);
      rematch006_in_bus_rdat_last  : in  std_logic;
      rematch006_in_cmd_valid      : in  std_logic;
      rematch006_in_cmd_ready      : out std_logic;
      rematch006_in_cmd_firstIdx   : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch006_in_cmd_lastIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch006_in_cmd_ctrl       : in  std_logic_vector(REMATCH006_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch006_in_cmd_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch006_in_unl_valid      : out std_logic;
      rematch006_in_unl_ready      : in  std_logic;
      rematch006_in_unl_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  component Kernel_rematch007 is
    generic (
      INDEX_WIDTH                      : integer := 32;
      TAG_WIDTH                        : integer := 1;
      REMATCH007_IN_BUS_ADDR_WIDTH     : integer := 64;
      REMATCH007_IN_BUS_DATA_WIDTH     : integer := 512;
      REMATCH007_IN_BUS_LEN_WIDTH      : integer := 8;
      REMATCH007_IN_BUS_BURST_STEP_LEN : integer := 1;
      REMATCH007_IN_BUS_BURST_MAX_LEN  : integer := 16
    );
    port (
      bcd_clk                      : in  std_logic;
      bcd_reset                    : in  std_logic;
      kcd_clk                      : in  std_logic;
      kcd_reset                    : in  std_logic;
      rematch007_in_valid          : out std_logic;
      rematch007_in_ready          : in  std_logic;
      rematch007_in_dvalid         : out std_logic;
      rematch007_in_last           : out std_logic;
      rematch007_in_length         : out std_logic_vector(31 downto 0);
      rematch007_in_count          : out std_logic_vector(0 downto 0);
      rematch007_in_chars_valid    : out std_logic;
      rematch007_in_chars_ready    : in  std_logic;
      rematch007_in_chars_dvalid   : out std_logic;
      rematch007_in_chars_last     : out std_logic;
      rematch007_in_chars          : out std_logic_vector(31 downto 0);
      rematch007_in_chars_count    : out std_logic_vector(2 downto 0);
      rematch007_in_bus_rreq_valid : out std_logic;
      rematch007_in_bus_rreq_ready : in  std_logic;
      rematch007_in_bus_rreq_addr  : out std_logic_vector(REMATCH007_IN_BUS_ADDR_WIDTH-1 downto 0);
      rematch007_in_bus_rreq_len   : out std_logic_vector(REMATCH007_IN_BUS_LEN_WIDTH-1 downto 0);
      rematch007_in_bus_rdat_valid : in  std_logic;
      rematch007_in_bus_rdat_ready : out std_logic;
      rematch007_in_bus_rdat_data  : in  std_logic_vector(REMATCH007_IN_BUS_DATA_WIDTH-1 downto 0);
      rematch007_in_bus_rdat_last  : in  std_logic;
      rematch007_in_cmd_valid      : in  std_logic;
      rematch007_in_cmd_ready      : out std_logic;
      rematch007_in_cmd_firstIdx   : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch007_in_cmd_lastIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch007_in_cmd_ctrl       : in  std_logic_vector(REMATCH007_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch007_in_cmd_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch007_in_unl_valid      : out std_logic;
      rematch007_in_unl_ready      : in  std_logic;
      rematch007_in_unl_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  component Kernel_rematch008 is
    generic (
      INDEX_WIDTH                      : integer := 32;
      TAG_WIDTH                        : integer := 1;
      REMATCH008_IN_BUS_ADDR_WIDTH     : integer := 64;
      REMATCH008_IN_BUS_DATA_WIDTH     : integer := 512;
      REMATCH008_IN_BUS_LEN_WIDTH      : integer := 8;
      REMATCH008_IN_BUS_BURST_STEP_LEN : integer := 1;
      REMATCH008_IN_BUS_BURST_MAX_LEN  : integer := 16
    );
    port (
      bcd_clk                      : in  std_logic;
      bcd_reset                    : in  std_logic;
      kcd_clk                      : in  std_logic;
      kcd_reset                    : in  std_logic;
      rematch008_in_valid          : out std_logic;
      rematch008_in_ready          : in  std_logic;
      rematch008_in_dvalid         : out std_logic;
      rematch008_in_last           : out std_logic;
      rematch008_in_length         : out std_logic_vector(31 downto 0);
      rematch008_in_count          : out std_logic_vector(0 downto 0);
      rematch008_in_chars_valid    : out std_logic;
      rematch008_in_chars_ready    : in  std_logic;
      rematch008_in_chars_dvalid   : out std_logic;
      rematch008_in_chars_last     : out std_logic;
      rematch008_in_chars          : out std_logic_vector(31 downto 0);
      rematch008_in_chars_count    : out std_logic_vector(2 downto 0);
      rematch008_in_bus_rreq_valid : out std_logic;
      rematch008_in_bus_rreq_ready : in  std_logic;
      rematch008_in_bus_rreq_addr  : out std_logic_vector(REMATCH008_IN_BUS_ADDR_WIDTH-1 downto 0);
      rematch008_in_bus_rreq_len   : out std_logic_vector(REMATCH008_IN_BUS_LEN_WIDTH-1 downto 0);
      rematch008_in_bus_rdat_valid : in  std_logic;
      rematch008_in_bus_rdat_ready : out std_logic;
      rematch008_in_bus_rdat_data  : in  std_logic_vector(REMATCH008_IN_BUS_DATA_WIDTH-1 downto 0);
      rematch008_in_bus_rdat_last  : in  std_logic;
      rematch008_in_cmd_valid      : in  std_logic;
      rematch008_in_cmd_ready      : out std_logic;
      rematch008_in_cmd_firstIdx   : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch008_in_cmd_lastIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch008_in_cmd_ctrl       : in  std_logic_vector(REMATCH008_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch008_in_cmd_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch008_in_unl_valid      : out std_logic;
      rematch008_in_unl_ready      : in  std_logic;
      rematch008_in_unl_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  component Kernel_rematch009 is
    generic (
      INDEX_WIDTH                      : integer := 32;
      TAG_WIDTH                        : integer := 1;
      REMATCH009_IN_BUS_ADDR_WIDTH     : integer := 64;
      REMATCH009_IN_BUS_DATA_WIDTH     : integer := 512;
      REMATCH009_IN_BUS_LEN_WIDTH      : integer := 8;
      REMATCH009_IN_BUS_BURST_STEP_LEN : integer := 1;
      REMATCH009_IN_BUS_BURST_MAX_LEN  : integer := 16
    );
    port (
      bcd_clk                      : in  std_logic;
      bcd_reset                    : in  std_logic;
      kcd_clk                      : in  std_logic;
      kcd_reset                    : in  std_logic;
      rematch009_in_valid          : out std_logic;
      rematch009_in_ready          : in  std_logic;
      rematch009_in_dvalid         : out std_logic;
      rematch009_in_last           : out std_logic;
      rematch009_in_length         : out std_logic_vector(31 downto 0);
      rematch009_in_count          : out std_logic_vector(0 downto 0);
      rematch009_in_chars_valid    : out std_logic;
      rematch009_in_chars_ready    : in  std_logic;
      rematch009_in_chars_dvalid   : out std_logic;
      rematch009_in_chars_last     : out std_logic;
      rematch009_in_chars          : out std_logic_vector(31 downto 0);
      rematch009_in_chars_count    : out std_logic_vector(2 downto 0);
      rematch009_in_bus_rreq_valid : out std_logic;
      rematch009_in_bus_rreq_ready : in  std_logic;
      rematch009_in_bus_rreq_addr  : out std_logic_vector(REMATCH009_IN_BUS_ADDR_WIDTH-1 downto 0);
      rematch009_in_bus_rreq_len   : out std_logic_vector(REMATCH009_IN_BUS_LEN_WIDTH-1 downto 0);
      rematch009_in_bus_rdat_valid : in  std_logic;
      rematch009_in_bus_rdat_ready : out std_logic;
      rematch009_in_bus_rdat_data  : in  std_logic_vector(REMATCH009_IN_BUS_DATA_WIDTH-1 downto 0);
      rematch009_in_bus_rdat_last  : in  std_logic;
      rematch009_in_cmd_valid      : in  std_logic;
      rematch009_in_cmd_ready      : out std_logic;
      rematch009_in_cmd_firstIdx   : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch009_in_cmd_lastIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch009_in_cmd_ctrl       : in  std_logic_vector(REMATCH009_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch009_in_cmd_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch009_in_unl_valid      : out std_logic;
      rematch009_in_unl_ready      : in  std_logic;
      rematch009_in_unl_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  component Kernel_rematch010 is
    generic (
      INDEX_WIDTH                      : integer := 32;
      TAG_WIDTH                        : integer := 1;
      REMATCH010_IN_BUS_ADDR_WIDTH     : integer := 64;
      REMATCH010_IN_BUS_DATA_WIDTH     : integer := 512;
      REMATCH010_IN_BUS_LEN_WIDTH      : integer := 8;
      REMATCH010_IN_BUS_BURST_STEP_LEN : integer := 1;
      REMATCH010_IN_BUS_BURST_MAX_LEN  : integer := 16
    );
    port (
      bcd_clk                      : in  std_logic;
      bcd_reset                    : in  std_logic;
      kcd_clk                      : in  std_logic;
      kcd_reset                    : in  std_logic;
      rematch010_in_valid          : out std_logic;
      rematch010_in_ready          : in  std_logic;
      rematch010_in_dvalid         : out std_logic;
      rematch010_in_last           : out std_logic;
      rematch010_in_length         : out std_logic_vector(31 downto 0);
      rematch010_in_count          : out std_logic_vector(0 downto 0);
      rematch010_in_chars_valid    : out std_logic;
      rematch010_in_chars_ready    : in  std_logic;
      rematch010_in_chars_dvalid   : out std_logic;
      rematch010_in_chars_last     : out std_logic;
      rematch010_in_chars          : out std_logic_vector(31 downto 0);
      rematch010_in_chars_count    : out std_logic_vector(2 downto 0);
      rematch010_in_bus_rreq_valid : out std_logic;
      rematch010_in_bus_rreq_ready : in  std_logic;
      rematch010_in_bus_rreq_addr  : out std_logic_vector(REMATCH010_IN_BUS_ADDR_WIDTH-1 downto 0);
      rematch010_in_bus_rreq_len   : out std_logic_vector(REMATCH010_IN_BUS_LEN_WIDTH-1 downto 0);
      rematch010_in_bus_rdat_valid : in  std_logic;
      rematch010_in_bus_rdat_ready : out std_logic;
      rematch010_in_bus_rdat_data  : in  std_logic_vector(REMATCH010_IN_BUS_DATA_WIDTH-1 downto 0);
      rematch010_in_bus_rdat_last  : in  std_logic;
      rematch010_in_cmd_valid      : in  std_logic;
      rematch010_in_cmd_ready      : out std_logic;
      rematch010_in_cmd_firstIdx   : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch010_in_cmd_lastIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch010_in_cmd_ctrl       : in  std_logic_vector(REMATCH010_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch010_in_cmd_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch010_in_unl_valid      : out std_logic;
      rematch010_in_unl_ready      : in  std_logic;
      rematch010_in_unl_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  component Kernel_rematch011 is
    generic (
      INDEX_WIDTH                      : integer := 32;
      TAG_WIDTH                        : integer := 1;
      REMATCH011_IN_BUS_ADDR_WIDTH     : integer := 64;
      REMATCH011_IN_BUS_DATA_WIDTH     : integer := 512;
      REMATCH011_IN_BUS_LEN_WIDTH      : integer := 8;
      REMATCH011_IN_BUS_BURST_STEP_LEN : integer := 1;
      REMATCH011_IN_BUS_BURST_MAX_LEN  : integer := 16
    );
    port (
      bcd_clk                      : in  std_logic;
      bcd_reset                    : in  std_logic;
      kcd_clk                      : in  std_logic;
      kcd_reset                    : in  std_logic;
      rematch011_in_valid          : out std_logic;
      rematch011_in_ready          : in  std_logic;
      rematch011_in_dvalid         : out std_logic;
      rematch011_in_last           : out std_logic;
      rematch011_in_length         : out std_logic_vector(31 downto 0);
      rematch011_in_count          : out std_logic_vector(0 downto 0);
      rematch011_in_chars_valid    : out std_logic;
      rematch011_in_chars_ready    : in  std_logic;
      rematch011_in_chars_dvalid   : out std_logic;
      rematch011_in_chars_last     : out std_logic;
      rematch011_in_chars          : out std_logic_vector(31 downto 0);
      rematch011_in_chars_count    : out std_logic_vector(2 downto 0);
      rematch011_in_bus_rreq_valid : out std_logic;
      rematch011_in_bus_rreq_ready : in  std_logic;
      rematch011_in_bus_rreq_addr  : out std_logic_vector(REMATCH011_IN_BUS_ADDR_WIDTH-1 downto 0);
      rematch011_in_bus_rreq_len   : out std_logic_vector(REMATCH011_IN_BUS_LEN_WIDTH-1 downto 0);
      rematch011_in_bus_rdat_valid : in  std_logic;
      rematch011_in_bus_rdat_ready : out std_logic;
      rematch011_in_bus_rdat_data  : in  std_logic_vector(REMATCH011_IN_BUS_DATA_WIDTH-1 downto 0);
      rematch011_in_bus_rdat_last  : in  std_logic;
      rematch011_in_cmd_valid      : in  std_logic;
      rematch011_in_cmd_ready      : out std_logic;
      rematch011_in_cmd_firstIdx   : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch011_in_cmd_lastIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch011_in_cmd_ctrl       : in  std_logic_vector(REMATCH011_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch011_in_cmd_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch011_in_unl_valid      : out std_logic;
      rematch011_in_unl_ready      : in  std_logic;
      rematch011_in_unl_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  component Kernel_rematch012 is
    generic (
      INDEX_WIDTH                      : integer := 32;
      TAG_WIDTH                        : integer := 1;
      REMATCH012_IN_BUS_ADDR_WIDTH     : integer := 64;
      REMATCH012_IN_BUS_DATA_WIDTH     : integer := 512;
      REMATCH012_IN_BUS_LEN_WIDTH      : integer := 8;
      REMATCH012_IN_BUS_BURST_STEP_LEN : integer := 1;
      REMATCH012_IN_BUS_BURST_MAX_LEN  : integer := 16
    );
    port (
      bcd_clk                      : in  std_logic;
      bcd_reset                    : in  std_logic;
      kcd_clk                      : in  std_logic;
      kcd_reset                    : in  std_logic;
      rematch012_in_valid          : out std_logic;
      rematch012_in_ready          : in  std_logic;
      rematch012_in_dvalid         : out std_logic;
      rematch012_in_last           : out std_logic;
      rematch012_in_length         : out std_logic_vector(31 downto 0);
      rematch012_in_count          : out std_logic_vector(0 downto 0);
      rematch012_in_chars_valid    : out std_logic;
      rematch012_in_chars_ready    : in  std_logic;
      rematch012_in_chars_dvalid   : out std_logic;
      rematch012_in_chars_last     : out std_logic;
      rematch012_in_chars          : out std_logic_vector(31 downto 0);
      rematch012_in_chars_count    : out std_logic_vector(2 downto 0);
      rematch012_in_bus_rreq_valid : out std_logic;
      rematch012_in_bus_rreq_ready : in  std_logic;
      rematch012_in_bus_rreq_addr  : out std_logic_vector(REMATCH012_IN_BUS_ADDR_WIDTH-1 downto 0);
      rematch012_in_bus_rreq_len   : out std_logic_vector(REMATCH012_IN_BUS_LEN_WIDTH-1 downto 0);
      rematch012_in_bus_rdat_valid : in  std_logic;
      rematch012_in_bus_rdat_ready : out std_logic;
      rematch012_in_bus_rdat_data  : in  std_logic_vector(REMATCH012_IN_BUS_DATA_WIDTH-1 downto 0);
      rematch012_in_bus_rdat_last  : in  std_logic;
      rematch012_in_cmd_valid      : in  std_logic;
      rematch012_in_cmd_ready      : out std_logic;
      rematch012_in_cmd_firstIdx   : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch012_in_cmd_lastIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch012_in_cmd_ctrl       : in  std_logic_vector(REMATCH012_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch012_in_cmd_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch012_in_unl_valid      : out std_logic;
      rematch012_in_unl_ready      : in  std_logic;
      rematch012_in_unl_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  component Kernel_rematch013 is
    generic (
      INDEX_WIDTH                      : integer := 32;
      TAG_WIDTH                        : integer := 1;
      REMATCH013_IN_BUS_ADDR_WIDTH     : integer := 64;
      REMATCH013_IN_BUS_DATA_WIDTH     : integer := 512;
      REMATCH013_IN_BUS_LEN_WIDTH      : integer := 8;
      REMATCH013_IN_BUS_BURST_STEP_LEN : integer := 1;
      REMATCH013_IN_BUS_BURST_MAX_LEN  : integer := 16
    );
    port (
      bcd_clk                      : in  std_logic;
      bcd_reset                    : in  std_logic;
      kcd_clk                      : in  std_logic;
      kcd_reset                    : in  std_logic;
      rematch013_in_valid          : out std_logic;
      rematch013_in_ready          : in  std_logic;
      rematch013_in_dvalid         : out std_logic;
      rematch013_in_last           : out std_logic;
      rematch013_in_length         : out std_logic_vector(31 downto 0);
      rematch013_in_count          : out std_logic_vector(0 downto 0);
      rematch013_in_chars_valid    : out std_logic;
      rematch013_in_chars_ready    : in  std_logic;
      rematch013_in_chars_dvalid   : out std_logic;
      rematch013_in_chars_last     : out std_logic;
      rematch013_in_chars          : out std_logic_vector(31 downto 0);
      rematch013_in_chars_count    : out std_logic_vector(2 downto 0);
      rematch013_in_bus_rreq_valid : out std_logic;
      rematch013_in_bus_rreq_ready : in  std_logic;
      rematch013_in_bus_rreq_addr  : out std_logic_vector(REMATCH013_IN_BUS_ADDR_WIDTH-1 downto 0);
      rematch013_in_bus_rreq_len   : out std_logic_vector(REMATCH013_IN_BUS_LEN_WIDTH-1 downto 0);
      rematch013_in_bus_rdat_valid : in  std_logic;
      rematch013_in_bus_rdat_ready : out std_logic;
      rematch013_in_bus_rdat_data  : in  std_logic_vector(REMATCH013_IN_BUS_DATA_WIDTH-1 downto 0);
      rematch013_in_bus_rdat_last  : in  std_logic;
      rematch013_in_cmd_valid      : in  std_logic;
      rematch013_in_cmd_ready      : out std_logic;
      rematch013_in_cmd_firstIdx   : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch013_in_cmd_lastIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch013_in_cmd_ctrl       : in  std_logic_vector(REMATCH013_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch013_in_cmd_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch013_in_unl_valid      : out std_logic;
      rematch013_in_unl_ready      : in  std_logic;
      rematch013_in_unl_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  component Kernel_rematch014 is
    generic (
      INDEX_WIDTH                      : integer := 32;
      TAG_WIDTH                        : integer := 1;
      REMATCH014_IN_BUS_ADDR_WIDTH     : integer := 64;
      REMATCH014_IN_BUS_DATA_WIDTH     : integer := 512;
      REMATCH014_IN_BUS_LEN_WIDTH      : integer := 8;
      REMATCH014_IN_BUS_BURST_STEP_LEN : integer := 1;
      REMATCH014_IN_BUS_BURST_MAX_LEN  : integer := 16
    );
    port (
      bcd_clk                      : in  std_logic;
      bcd_reset                    : in  std_logic;
      kcd_clk                      : in  std_logic;
      kcd_reset                    : in  std_logic;
      rematch014_in_valid          : out std_logic;
      rematch014_in_ready          : in  std_logic;
      rematch014_in_dvalid         : out std_logic;
      rematch014_in_last           : out std_logic;
      rematch014_in_length         : out std_logic_vector(31 downto 0);
      rematch014_in_count          : out std_logic_vector(0 downto 0);
      rematch014_in_chars_valid    : out std_logic;
      rematch014_in_chars_ready    : in  std_logic;
      rematch014_in_chars_dvalid   : out std_logic;
      rematch014_in_chars_last     : out std_logic;
      rematch014_in_chars          : out std_logic_vector(31 downto 0);
      rematch014_in_chars_count    : out std_logic_vector(2 downto 0);
      rematch014_in_bus_rreq_valid : out std_logic;
      rematch014_in_bus_rreq_ready : in  std_logic;
      rematch014_in_bus_rreq_addr  : out std_logic_vector(REMATCH014_IN_BUS_ADDR_WIDTH-1 downto 0);
      rematch014_in_bus_rreq_len   : out std_logic_vector(REMATCH014_IN_BUS_LEN_WIDTH-1 downto 0);
      rematch014_in_bus_rdat_valid : in  std_logic;
      rematch014_in_bus_rdat_ready : out std_logic;
      rematch014_in_bus_rdat_data  : in  std_logic_vector(REMATCH014_IN_BUS_DATA_WIDTH-1 downto 0);
      rematch014_in_bus_rdat_last  : in  std_logic;
      rematch014_in_cmd_valid      : in  std_logic;
      rematch014_in_cmd_ready      : out std_logic;
      rematch014_in_cmd_firstIdx   : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch014_in_cmd_lastIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch014_in_cmd_ctrl       : in  std_logic_vector(REMATCH014_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch014_in_cmd_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch014_in_unl_valid      : out std_logic;
      rematch014_in_unl_ready      : in  std_logic;
      rematch014_in_unl_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  component Kernel_rematch015 is
    generic (
      INDEX_WIDTH                      : integer := 32;
      TAG_WIDTH                        : integer := 1;
      REMATCH015_IN_BUS_ADDR_WIDTH     : integer := 64;
      REMATCH015_IN_BUS_DATA_WIDTH     : integer := 512;
      REMATCH015_IN_BUS_LEN_WIDTH      : integer := 8;
      REMATCH015_IN_BUS_BURST_STEP_LEN : integer := 1;
      REMATCH015_IN_BUS_BURST_MAX_LEN  : integer := 16
    );
    port (
      bcd_clk                      : in  std_logic;
      bcd_reset                    : in  std_logic;
      kcd_clk                      : in  std_logic;
      kcd_reset                    : in  std_logic;
      rematch015_in_valid          : out std_logic;
      rematch015_in_ready          : in  std_logic;
      rematch015_in_dvalid         : out std_logic;
      rematch015_in_last           : out std_logic;
      rematch015_in_length         : out std_logic_vector(31 downto 0);
      rematch015_in_count          : out std_logic_vector(0 downto 0);
      rematch015_in_chars_valid    : out std_logic;
      rematch015_in_chars_ready    : in  std_logic;
      rematch015_in_chars_dvalid   : out std_logic;
      rematch015_in_chars_last     : out std_logic;
      rematch015_in_chars          : out std_logic_vector(31 downto 0);
      rematch015_in_chars_count    : out std_logic_vector(2 downto 0);
      rematch015_in_bus_rreq_valid : out std_logic;
      rematch015_in_bus_rreq_ready : in  std_logic;
      rematch015_in_bus_rreq_addr  : out std_logic_vector(REMATCH015_IN_BUS_ADDR_WIDTH-1 downto 0);
      rematch015_in_bus_rreq_len   : out std_logic_vector(REMATCH015_IN_BUS_LEN_WIDTH-1 downto 0);
      rematch015_in_bus_rdat_valid : in  std_logic;
      rematch015_in_bus_rdat_ready : out std_logic;
      rematch015_in_bus_rdat_data  : in  std_logic_vector(REMATCH015_IN_BUS_DATA_WIDTH-1 downto 0);
      rematch015_in_bus_rdat_last  : in  std_logic;
      rematch015_in_cmd_valid      : in  std_logic;
      rematch015_in_cmd_ready      : out std_logic;
      rematch015_in_cmd_firstIdx   : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch015_in_cmd_lastIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      rematch015_in_cmd_ctrl       : in  std_logic_vector(REMATCH015_IN_BUS_ADDR_WIDTH*2-1 downto 0);
      rematch015_in_cmd_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      rematch015_in_unl_valid      : out std_logic;
      rematch015_in_unl_ready      : in  std_logic;
      rematch015_in_unl_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  signal Kernel_Nucleus_inst_mmio_awvalid                    : std_logic;
  signal Kernel_Nucleus_inst_mmio_awready                    : std_logic;
  signal Kernel_Nucleus_inst_mmio_awaddr                     : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_mmio_wvalid                     : std_logic;
  signal Kernel_Nucleus_inst_mmio_wready                     : std_logic;
  signal Kernel_Nucleus_inst_mmio_wdata                      : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_mmio_wstrb                      : std_logic_vector(3 downto 0);
  signal Kernel_Nucleus_inst_mmio_bvalid                     : std_logic;
  signal Kernel_Nucleus_inst_mmio_bready                     : std_logic;
  signal Kernel_Nucleus_inst_mmio_bresp                      : std_logic_vector(1 downto 0);
  signal Kernel_Nucleus_inst_mmio_arvalid                    : std_logic;
  signal Kernel_Nucleus_inst_mmio_arready                    : std_logic;
  signal Kernel_Nucleus_inst_mmio_araddr                     : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_mmio_rvalid                     : std_logic;
  signal Kernel_Nucleus_inst_mmio_rready                     : std_logic;
  signal Kernel_Nucleus_inst_mmio_rdata                      : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_mmio_rresp                      : std_logic_vector(1 downto 0);

  signal Kernel_Nucleus_inst_rematch000_in_valid             : std_logic;
  signal Kernel_Nucleus_inst_rematch000_in_ready             : std_logic;
  signal Kernel_Nucleus_inst_rematch000_in_dvalid            : std_logic;
  signal Kernel_Nucleus_inst_rematch000_in_last              : std_logic;
  signal Kernel_Nucleus_inst_rematch000_in_length            : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch000_in_count             : std_logic_vector(0 downto 0);
  signal Kernel_Nucleus_inst_rematch000_in_chars_valid       : std_logic;
  signal Kernel_Nucleus_inst_rematch000_in_chars_ready       : std_logic;
  signal Kernel_Nucleus_inst_rematch000_in_chars_dvalid      : std_logic;
  signal Kernel_Nucleus_inst_rematch000_in_chars_last        : std_logic;
  signal Kernel_Nucleus_inst_rematch000_in_chars             : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch000_in_chars_count       : std_logic_vector(2 downto 0);

  signal Kernel_Nucleus_inst_rematch000_in_unl_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch000_in_unl_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch000_in_unl_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch000_in_cmd_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch000_in_cmd_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch000_in_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch000_in_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch000_in_cmd_ctrl          : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_Nucleus_inst_rematch000_in_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch001_in_valid             : std_logic;
  signal Kernel_Nucleus_inst_rematch001_in_ready             : std_logic;
  signal Kernel_Nucleus_inst_rematch001_in_dvalid            : std_logic;
  signal Kernel_Nucleus_inst_rematch001_in_last              : std_logic;
  signal Kernel_Nucleus_inst_rematch001_in_length            : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch001_in_count             : std_logic_vector(0 downto 0);
  signal Kernel_Nucleus_inst_rematch001_in_chars_valid       : std_logic;
  signal Kernel_Nucleus_inst_rematch001_in_chars_ready       : std_logic;
  signal Kernel_Nucleus_inst_rematch001_in_chars_dvalid      : std_logic;
  signal Kernel_Nucleus_inst_rematch001_in_chars_last        : std_logic;
  signal Kernel_Nucleus_inst_rematch001_in_chars             : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch001_in_chars_count       : std_logic_vector(2 downto 0);

  signal Kernel_Nucleus_inst_rematch001_in_unl_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch001_in_unl_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch001_in_unl_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch001_in_cmd_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch001_in_cmd_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch001_in_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch001_in_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch001_in_cmd_ctrl          : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_Nucleus_inst_rematch001_in_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch002_in_valid             : std_logic;
  signal Kernel_Nucleus_inst_rematch002_in_ready             : std_logic;
  signal Kernel_Nucleus_inst_rematch002_in_dvalid            : std_logic;
  signal Kernel_Nucleus_inst_rematch002_in_last              : std_logic;
  signal Kernel_Nucleus_inst_rematch002_in_length            : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch002_in_count             : std_logic_vector(0 downto 0);
  signal Kernel_Nucleus_inst_rematch002_in_chars_valid       : std_logic;
  signal Kernel_Nucleus_inst_rematch002_in_chars_ready       : std_logic;
  signal Kernel_Nucleus_inst_rematch002_in_chars_dvalid      : std_logic;
  signal Kernel_Nucleus_inst_rematch002_in_chars_last        : std_logic;
  signal Kernel_Nucleus_inst_rematch002_in_chars             : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch002_in_chars_count       : std_logic_vector(2 downto 0);

  signal Kernel_Nucleus_inst_rematch002_in_unl_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch002_in_unl_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch002_in_unl_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch002_in_cmd_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch002_in_cmd_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch002_in_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch002_in_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch002_in_cmd_ctrl          : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_Nucleus_inst_rematch002_in_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch003_in_valid             : std_logic;
  signal Kernel_Nucleus_inst_rematch003_in_ready             : std_logic;
  signal Kernel_Nucleus_inst_rematch003_in_dvalid            : std_logic;
  signal Kernel_Nucleus_inst_rematch003_in_last              : std_logic;
  signal Kernel_Nucleus_inst_rematch003_in_length            : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch003_in_count             : std_logic_vector(0 downto 0);
  signal Kernel_Nucleus_inst_rematch003_in_chars_valid       : std_logic;
  signal Kernel_Nucleus_inst_rematch003_in_chars_ready       : std_logic;
  signal Kernel_Nucleus_inst_rematch003_in_chars_dvalid      : std_logic;
  signal Kernel_Nucleus_inst_rematch003_in_chars_last        : std_logic;
  signal Kernel_Nucleus_inst_rematch003_in_chars             : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch003_in_chars_count       : std_logic_vector(2 downto 0);

  signal Kernel_Nucleus_inst_rematch003_in_unl_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch003_in_unl_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch003_in_unl_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch003_in_cmd_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch003_in_cmd_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch003_in_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch003_in_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch003_in_cmd_ctrl          : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_Nucleus_inst_rematch003_in_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch004_in_valid             : std_logic;
  signal Kernel_Nucleus_inst_rematch004_in_ready             : std_logic;
  signal Kernel_Nucleus_inst_rematch004_in_dvalid            : std_logic;
  signal Kernel_Nucleus_inst_rematch004_in_last              : std_logic;
  signal Kernel_Nucleus_inst_rematch004_in_length            : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch004_in_count             : std_logic_vector(0 downto 0);
  signal Kernel_Nucleus_inst_rematch004_in_chars_valid       : std_logic;
  signal Kernel_Nucleus_inst_rematch004_in_chars_ready       : std_logic;
  signal Kernel_Nucleus_inst_rematch004_in_chars_dvalid      : std_logic;
  signal Kernel_Nucleus_inst_rematch004_in_chars_last        : std_logic;
  signal Kernel_Nucleus_inst_rematch004_in_chars             : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch004_in_chars_count       : std_logic_vector(2 downto 0);

  signal Kernel_Nucleus_inst_rematch004_in_unl_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch004_in_unl_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch004_in_unl_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch004_in_cmd_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch004_in_cmd_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch004_in_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch004_in_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch004_in_cmd_ctrl          : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_Nucleus_inst_rematch004_in_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch005_in_valid             : std_logic;
  signal Kernel_Nucleus_inst_rematch005_in_ready             : std_logic;
  signal Kernel_Nucleus_inst_rematch005_in_dvalid            : std_logic;
  signal Kernel_Nucleus_inst_rematch005_in_last              : std_logic;
  signal Kernel_Nucleus_inst_rematch005_in_length            : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch005_in_count             : std_logic_vector(0 downto 0);
  signal Kernel_Nucleus_inst_rematch005_in_chars_valid       : std_logic;
  signal Kernel_Nucleus_inst_rematch005_in_chars_ready       : std_logic;
  signal Kernel_Nucleus_inst_rematch005_in_chars_dvalid      : std_logic;
  signal Kernel_Nucleus_inst_rematch005_in_chars_last        : std_logic;
  signal Kernel_Nucleus_inst_rematch005_in_chars             : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch005_in_chars_count       : std_logic_vector(2 downto 0);

  signal Kernel_Nucleus_inst_rematch005_in_unl_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch005_in_unl_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch005_in_unl_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch005_in_cmd_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch005_in_cmd_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch005_in_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch005_in_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch005_in_cmd_ctrl          : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_Nucleus_inst_rematch005_in_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch006_in_valid             : std_logic;
  signal Kernel_Nucleus_inst_rematch006_in_ready             : std_logic;
  signal Kernel_Nucleus_inst_rematch006_in_dvalid            : std_logic;
  signal Kernel_Nucleus_inst_rematch006_in_last              : std_logic;
  signal Kernel_Nucleus_inst_rematch006_in_length            : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch006_in_count             : std_logic_vector(0 downto 0);
  signal Kernel_Nucleus_inst_rematch006_in_chars_valid       : std_logic;
  signal Kernel_Nucleus_inst_rematch006_in_chars_ready       : std_logic;
  signal Kernel_Nucleus_inst_rematch006_in_chars_dvalid      : std_logic;
  signal Kernel_Nucleus_inst_rematch006_in_chars_last        : std_logic;
  signal Kernel_Nucleus_inst_rematch006_in_chars             : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch006_in_chars_count       : std_logic_vector(2 downto 0);

  signal Kernel_Nucleus_inst_rematch006_in_unl_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch006_in_unl_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch006_in_unl_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch006_in_cmd_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch006_in_cmd_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch006_in_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch006_in_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch006_in_cmd_ctrl          : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_Nucleus_inst_rematch006_in_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch007_in_valid             : std_logic;
  signal Kernel_Nucleus_inst_rematch007_in_ready             : std_logic;
  signal Kernel_Nucleus_inst_rematch007_in_dvalid            : std_logic;
  signal Kernel_Nucleus_inst_rematch007_in_last              : std_logic;
  signal Kernel_Nucleus_inst_rematch007_in_length            : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch007_in_count             : std_logic_vector(0 downto 0);
  signal Kernel_Nucleus_inst_rematch007_in_chars_valid       : std_logic;
  signal Kernel_Nucleus_inst_rematch007_in_chars_ready       : std_logic;
  signal Kernel_Nucleus_inst_rematch007_in_chars_dvalid      : std_logic;
  signal Kernel_Nucleus_inst_rematch007_in_chars_last        : std_logic;
  signal Kernel_Nucleus_inst_rematch007_in_chars             : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch007_in_chars_count       : std_logic_vector(2 downto 0);

  signal Kernel_Nucleus_inst_rematch007_in_unl_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch007_in_unl_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch007_in_unl_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch007_in_cmd_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch007_in_cmd_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch007_in_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch007_in_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch007_in_cmd_ctrl          : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_Nucleus_inst_rematch007_in_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch008_in_valid             : std_logic;
  signal Kernel_Nucleus_inst_rematch008_in_ready             : std_logic;
  signal Kernel_Nucleus_inst_rematch008_in_dvalid            : std_logic;
  signal Kernel_Nucleus_inst_rematch008_in_last              : std_logic;
  signal Kernel_Nucleus_inst_rematch008_in_length            : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch008_in_count             : std_logic_vector(0 downto 0);
  signal Kernel_Nucleus_inst_rematch008_in_chars_valid       : std_logic;
  signal Kernel_Nucleus_inst_rematch008_in_chars_ready       : std_logic;
  signal Kernel_Nucleus_inst_rematch008_in_chars_dvalid      : std_logic;
  signal Kernel_Nucleus_inst_rematch008_in_chars_last        : std_logic;
  signal Kernel_Nucleus_inst_rematch008_in_chars             : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch008_in_chars_count       : std_logic_vector(2 downto 0);

  signal Kernel_Nucleus_inst_rematch008_in_unl_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch008_in_unl_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch008_in_unl_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch008_in_cmd_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch008_in_cmd_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch008_in_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch008_in_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch008_in_cmd_ctrl          : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_Nucleus_inst_rematch008_in_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch009_in_valid             : std_logic;
  signal Kernel_Nucleus_inst_rematch009_in_ready             : std_logic;
  signal Kernel_Nucleus_inst_rematch009_in_dvalid            : std_logic;
  signal Kernel_Nucleus_inst_rematch009_in_last              : std_logic;
  signal Kernel_Nucleus_inst_rematch009_in_length            : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch009_in_count             : std_logic_vector(0 downto 0);
  signal Kernel_Nucleus_inst_rematch009_in_chars_valid       : std_logic;
  signal Kernel_Nucleus_inst_rematch009_in_chars_ready       : std_logic;
  signal Kernel_Nucleus_inst_rematch009_in_chars_dvalid      : std_logic;
  signal Kernel_Nucleus_inst_rematch009_in_chars_last        : std_logic;
  signal Kernel_Nucleus_inst_rematch009_in_chars             : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch009_in_chars_count       : std_logic_vector(2 downto 0);

  signal Kernel_Nucleus_inst_rematch009_in_unl_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch009_in_unl_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch009_in_unl_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch009_in_cmd_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch009_in_cmd_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch009_in_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch009_in_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch009_in_cmd_ctrl          : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_Nucleus_inst_rematch009_in_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch010_in_valid             : std_logic;
  signal Kernel_Nucleus_inst_rematch010_in_ready             : std_logic;
  signal Kernel_Nucleus_inst_rematch010_in_dvalid            : std_logic;
  signal Kernel_Nucleus_inst_rematch010_in_last              : std_logic;
  signal Kernel_Nucleus_inst_rematch010_in_length            : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch010_in_count             : std_logic_vector(0 downto 0);
  signal Kernel_Nucleus_inst_rematch010_in_chars_valid       : std_logic;
  signal Kernel_Nucleus_inst_rematch010_in_chars_ready       : std_logic;
  signal Kernel_Nucleus_inst_rematch010_in_chars_dvalid      : std_logic;
  signal Kernel_Nucleus_inst_rematch010_in_chars_last        : std_logic;
  signal Kernel_Nucleus_inst_rematch010_in_chars             : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch010_in_chars_count       : std_logic_vector(2 downto 0);

  signal Kernel_Nucleus_inst_rematch010_in_unl_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch010_in_unl_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch010_in_unl_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch010_in_cmd_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch010_in_cmd_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch010_in_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch010_in_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch010_in_cmd_ctrl          : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_Nucleus_inst_rematch010_in_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch011_in_valid             : std_logic;
  signal Kernel_Nucleus_inst_rematch011_in_ready             : std_logic;
  signal Kernel_Nucleus_inst_rematch011_in_dvalid            : std_logic;
  signal Kernel_Nucleus_inst_rematch011_in_last              : std_logic;
  signal Kernel_Nucleus_inst_rematch011_in_length            : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch011_in_count             : std_logic_vector(0 downto 0);
  signal Kernel_Nucleus_inst_rematch011_in_chars_valid       : std_logic;
  signal Kernel_Nucleus_inst_rematch011_in_chars_ready       : std_logic;
  signal Kernel_Nucleus_inst_rematch011_in_chars_dvalid      : std_logic;
  signal Kernel_Nucleus_inst_rematch011_in_chars_last        : std_logic;
  signal Kernel_Nucleus_inst_rematch011_in_chars             : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch011_in_chars_count       : std_logic_vector(2 downto 0);

  signal Kernel_Nucleus_inst_rematch011_in_unl_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch011_in_unl_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch011_in_unl_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch011_in_cmd_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch011_in_cmd_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch011_in_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch011_in_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch011_in_cmd_ctrl          : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_Nucleus_inst_rematch011_in_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch012_in_valid             : std_logic;
  signal Kernel_Nucleus_inst_rematch012_in_ready             : std_logic;
  signal Kernel_Nucleus_inst_rematch012_in_dvalid            : std_logic;
  signal Kernel_Nucleus_inst_rematch012_in_last              : std_logic;
  signal Kernel_Nucleus_inst_rematch012_in_length            : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch012_in_count             : std_logic_vector(0 downto 0);
  signal Kernel_Nucleus_inst_rematch012_in_chars_valid       : std_logic;
  signal Kernel_Nucleus_inst_rematch012_in_chars_ready       : std_logic;
  signal Kernel_Nucleus_inst_rematch012_in_chars_dvalid      : std_logic;
  signal Kernel_Nucleus_inst_rematch012_in_chars_last        : std_logic;
  signal Kernel_Nucleus_inst_rematch012_in_chars             : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch012_in_chars_count       : std_logic_vector(2 downto 0);

  signal Kernel_Nucleus_inst_rematch012_in_unl_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch012_in_unl_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch012_in_unl_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch012_in_cmd_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch012_in_cmd_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch012_in_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch012_in_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch012_in_cmd_ctrl          : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_Nucleus_inst_rematch012_in_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch013_in_valid             : std_logic;
  signal Kernel_Nucleus_inst_rematch013_in_ready             : std_logic;
  signal Kernel_Nucleus_inst_rematch013_in_dvalid            : std_logic;
  signal Kernel_Nucleus_inst_rematch013_in_last              : std_logic;
  signal Kernel_Nucleus_inst_rematch013_in_length            : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch013_in_count             : std_logic_vector(0 downto 0);
  signal Kernel_Nucleus_inst_rematch013_in_chars_valid       : std_logic;
  signal Kernel_Nucleus_inst_rematch013_in_chars_ready       : std_logic;
  signal Kernel_Nucleus_inst_rematch013_in_chars_dvalid      : std_logic;
  signal Kernel_Nucleus_inst_rematch013_in_chars_last        : std_logic;
  signal Kernel_Nucleus_inst_rematch013_in_chars             : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch013_in_chars_count       : std_logic_vector(2 downto 0);

  signal Kernel_Nucleus_inst_rematch013_in_unl_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch013_in_unl_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch013_in_unl_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch013_in_cmd_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch013_in_cmd_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch013_in_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch013_in_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch013_in_cmd_ctrl          : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_Nucleus_inst_rematch013_in_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch014_in_valid             : std_logic;
  signal Kernel_Nucleus_inst_rematch014_in_ready             : std_logic;
  signal Kernel_Nucleus_inst_rematch014_in_dvalid            : std_logic;
  signal Kernel_Nucleus_inst_rematch014_in_last              : std_logic;
  signal Kernel_Nucleus_inst_rematch014_in_length            : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch014_in_count             : std_logic_vector(0 downto 0);
  signal Kernel_Nucleus_inst_rematch014_in_chars_valid       : std_logic;
  signal Kernel_Nucleus_inst_rematch014_in_chars_ready       : std_logic;
  signal Kernel_Nucleus_inst_rematch014_in_chars_dvalid      : std_logic;
  signal Kernel_Nucleus_inst_rematch014_in_chars_last        : std_logic;
  signal Kernel_Nucleus_inst_rematch014_in_chars             : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch014_in_chars_count       : std_logic_vector(2 downto 0);

  signal Kernel_Nucleus_inst_rematch014_in_unl_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch014_in_unl_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch014_in_unl_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch014_in_cmd_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch014_in_cmd_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch014_in_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch014_in_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch014_in_cmd_ctrl          : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_Nucleus_inst_rematch014_in_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch015_in_valid             : std_logic;
  signal Kernel_Nucleus_inst_rematch015_in_ready             : std_logic;
  signal Kernel_Nucleus_inst_rematch015_in_dvalid            : std_logic;
  signal Kernel_Nucleus_inst_rematch015_in_last              : std_logic;
  signal Kernel_Nucleus_inst_rematch015_in_length            : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch015_in_count             : std_logic_vector(0 downto 0);
  signal Kernel_Nucleus_inst_rematch015_in_chars_valid       : std_logic;
  signal Kernel_Nucleus_inst_rematch015_in_chars_ready       : std_logic;
  signal Kernel_Nucleus_inst_rematch015_in_chars_dvalid      : std_logic;
  signal Kernel_Nucleus_inst_rematch015_in_chars_last        : std_logic;
  signal Kernel_Nucleus_inst_rematch015_in_chars             : std_logic_vector(31 downto 0);
  signal Kernel_Nucleus_inst_rematch015_in_chars_count       : std_logic_vector(2 downto 0);

  signal Kernel_Nucleus_inst_rematch015_in_unl_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch015_in_unl_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch015_in_unl_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_Nucleus_inst_rematch015_in_cmd_valid         : std_logic;
  signal Kernel_Nucleus_inst_rematch015_in_cmd_ready         : std_logic;
  signal Kernel_Nucleus_inst_rematch015_in_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch015_in_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_Nucleus_inst_rematch015_in_cmd_ctrl          : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_Nucleus_inst_rematch015_in_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch000_inst_rematch000_in_valid          : std_logic;
  signal Kernel_rematch000_inst_rematch000_in_ready          : std_logic;
  signal Kernel_rematch000_inst_rematch000_in_dvalid         : std_logic;
  signal Kernel_rematch000_inst_rematch000_in_last           : std_logic;
  signal Kernel_rematch000_inst_rematch000_in_length         : std_logic_vector(31 downto 0);
  signal Kernel_rematch000_inst_rematch000_in_count          : std_logic_vector(0 downto 0);
  signal Kernel_rematch000_inst_rematch000_in_chars_valid    : std_logic;
  signal Kernel_rematch000_inst_rematch000_in_chars_ready    : std_logic;
  signal Kernel_rematch000_inst_rematch000_in_chars_dvalid   : std_logic;
  signal Kernel_rematch000_inst_rematch000_in_chars_last     : std_logic;
  signal Kernel_rematch000_inst_rematch000_in_chars          : std_logic_vector(31 downto 0);
  signal Kernel_rematch000_inst_rematch000_in_chars_count    : std_logic_vector(2 downto 0);

  signal Kernel_rematch000_inst_rematch000_in_bus_rreq_valid : std_logic;
  signal Kernel_rematch000_inst_rematch000_in_bus_rreq_ready : std_logic;
  signal Kernel_rematch000_inst_rematch000_in_bus_rreq_addr  : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Kernel_rematch000_inst_rematch000_in_bus_rreq_len   : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Kernel_rematch000_inst_rematch000_in_bus_rdat_valid : std_logic;
  signal Kernel_rematch000_inst_rematch000_in_bus_rdat_ready : std_logic;
  signal Kernel_rematch000_inst_rematch000_in_bus_rdat_data  : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Kernel_rematch000_inst_rematch000_in_bus_rdat_last  : std_logic;

  signal Kernel_rematch000_inst_rematch000_in_cmd_valid      : std_logic;
  signal Kernel_rematch000_inst_rematch000_in_cmd_ready      : std_logic;
  signal Kernel_rematch000_inst_rematch000_in_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch000_inst_rematch000_in_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch000_inst_rematch000_in_cmd_ctrl       : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_rematch000_inst_rematch000_in_cmd_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch000_inst_rematch000_in_unl_valid      : std_logic;
  signal Kernel_rematch000_inst_rematch000_in_unl_ready      : std_logic;
  signal Kernel_rematch000_inst_rematch000_in_unl_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch001_inst_rematch001_in_valid          : std_logic;
  signal Kernel_rematch001_inst_rematch001_in_ready          : std_logic;
  signal Kernel_rematch001_inst_rematch001_in_dvalid         : std_logic;
  signal Kernel_rematch001_inst_rematch001_in_last           : std_logic;
  signal Kernel_rematch001_inst_rematch001_in_length         : std_logic_vector(31 downto 0);
  signal Kernel_rematch001_inst_rematch001_in_count          : std_logic_vector(0 downto 0);
  signal Kernel_rematch001_inst_rematch001_in_chars_valid    : std_logic;
  signal Kernel_rematch001_inst_rematch001_in_chars_ready    : std_logic;
  signal Kernel_rematch001_inst_rematch001_in_chars_dvalid   : std_logic;
  signal Kernel_rematch001_inst_rematch001_in_chars_last     : std_logic;
  signal Kernel_rematch001_inst_rematch001_in_chars          : std_logic_vector(31 downto 0);
  signal Kernel_rematch001_inst_rematch001_in_chars_count    : std_logic_vector(2 downto 0);

  signal Kernel_rematch001_inst_rematch001_in_bus_rreq_valid : std_logic;
  signal Kernel_rematch001_inst_rematch001_in_bus_rreq_ready : std_logic;
  signal Kernel_rematch001_inst_rematch001_in_bus_rreq_addr  : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Kernel_rematch001_inst_rematch001_in_bus_rreq_len   : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Kernel_rematch001_inst_rematch001_in_bus_rdat_valid : std_logic;
  signal Kernel_rematch001_inst_rematch001_in_bus_rdat_ready : std_logic;
  signal Kernel_rematch001_inst_rematch001_in_bus_rdat_data  : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Kernel_rematch001_inst_rematch001_in_bus_rdat_last  : std_logic;

  signal Kernel_rematch001_inst_rematch001_in_cmd_valid      : std_logic;
  signal Kernel_rematch001_inst_rematch001_in_cmd_ready      : std_logic;
  signal Kernel_rematch001_inst_rematch001_in_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch001_inst_rematch001_in_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch001_inst_rematch001_in_cmd_ctrl       : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_rematch001_inst_rematch001_in_cmd_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch001_inst_rematch001_in_unl_valid      : std_logic;
  signal Kernel_rematch001_inst_rematch001_in_unl_ready      : std_logic;
  signal Kernel_rematch001_inst_rematch001_in_unl_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch002_inst_rematch002_in_valid          : std_logic;
  signal Kernel_rematch002_inst_rematch002_in_ready          : std_logic;
  signal Kernel_rematch002_inst_rematch002_in_dvalid         : std_logic;
  signal Kernel_rematch002_inst_rematch002_in_last           : std_logic;
  signal Kernel_rematch002_inst_rematch002_in_length         : std_logic_vector(31 downto 0);
  signal Kernel_rematch002_inst_rematch002_in_count          : std_logic_vector(0 downto 0);
  signal Kernel_rematch002_inst_rematch002_in_chars_valid    : std_logic;
  signal Kernel_rematch002_inst_rematch002_in_chars_ready    : std_logic;
  signal Kernel_rematch002_inst_rematch002_in_chars_dvalid   : std_logic;
  signal Kernel_rematch002_inst_rematch002_in_chars_last     : std_logic;
  signal Kernel_rematch002_inst_rematch002_in_chars          : std_logic_vector(31 downto 0);
  signal Kernel_rematch002_inst_rematch002_in_chars_count    : std_logic_vector(2 downto 0);

  signal Kernel_rematch002_inst_rematch002_in_bus_rreq_valid : std_logic;
  signal Kernel_rematch002_inst_rematch002_in_bus_rreq_ready : std_logic;
  signal Kernel_rematch002_inst_rematch002_in_bus_rreq_addr  : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Kernel_rematch002_inst_rematch002_in_bus_rreq_len   : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Kernel_rematch002_inst_rematch002_in_bus_rdat_valid : std_logic;
  signal Kernel_rematch002_inst_rematch002_in_bus_rdat_ready : std_logic;
  signal Kernel_rematch002_inst_rematch002_in_bus_rdat_data  : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Kernel_rematch002_inst_rematch002_in_bus_rdat_last  : std_logic;

  signal Kernel_rematch002_inst_rematch002_in_cmd_valid      : std_logic;
  signal Kernel_rematch002_inst_rematch002_in_cmd_ready      : std_logic;
  signal Kernel_rematch002_inst_rematch002_in_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch002_inst_rematch002_in_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch002_inst_rematch002_in_cmd_ctrl       : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_rematch002_inst_rematch002_in_cmd_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch002_inst_rematch002_in_unl_valid      : std_logic;
  signal Kernel_rematch002_inst_rematch002_in_unl_ready      : std_logic;
  signal Kernel_rematch002_inst_rematch002_in_unl_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch003_inst_rematch003_in_valid          : std_logic;
  signal Kernel_rematch003_inst_rematch003_in_ready          : std_logic;
  signal Kernel_rematch003_inst_rematch003_in_dvalid         : std_logic;
  signal Kernel_rematch003_inst_rematch003_in_last           : std_logic;
  signal Kernel_rematch003_inst_rematch003_in_length         : std_logic_vector(31 downto 0);
  signal Kernel_rematch003_inst_rematch003_in_count          : std_logic_vector(0 downto 0);
  signal Kernel_rematch003_inst_rematch003_in_chars_valid    : std_logic;
  signal Kernel_rematch003_inst_rematch003_in_chars_ready    : std_logic;
  signal Kernel_rematch003_inst_rematch003_in_chars_dvalid   : std_logic;
  signal Kernel_rematch003_inst_rematch003_in_chars_last     : std_logic;
  signal Kernel_rematch003_inst_rematch003_in_chars          : std_logic_vector(31 downto 0);
  signal Kernel_rematch003_inst_rematch003_in_chars_count    : std_logic_vector(2 downto 0);

  signal Kernel_rematch003_inst_rematch003_in_bus_rreq_valid : std_logic;
  signal Kernel_rematch003_inst_rematch003_in_bus_rreq_ready : std_logic;
  signal Kernel_rematch003_inst_rematch003_in_bus_rreq_addr  : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Kernel_rematch003_inst_rematch003_in_bus_rreq_len   : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Kernel_rematch003_inst_rematch003_in_bus_rdat_valid : std_logic;
  signal Kernel_rematch003_inst_rematch003_in_bus_rdat_ready : std_logic;
  signal Kernel_rematch003_inst_rematch003_in_bus_rdat_data  : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Kernel_rematch003_inst_rematch003_in_bus_rdat_last  : std_logic;

  signal Kernel_rematch003_inst_rematch003_in_cmd_valid      : std_logic;
  signal Kernel_rematch003_inst_rematch003_in_cmd_ready      : std_logic;
  signal Kernel_rematch003_inst_rematch003_in_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch003_inst_rematch003_in_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch003_inst_rematch003_in_cmd_ctrl       : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_rematch003_inst_rematch003_in_cmd_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch003_inst_rematch003_in_unl_valid      : std_logic;
  signal Kernel_rematch003_inst_rematch003_in_unl_ready      : std_logic;
  signal Kernel_rematch003_inst_rematch003_in_unl_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch004_inst_rematch004_in_valid          : std_logic;
  signal Kernel_rematch004_inst_rematch004_in_ready          : std_logic;
  signal Kernel_rematch004_inst_rematch004_in_dvalid         : std_logic;
  signal Kernel_rematch004_inst_rematch004_in_last           : std_logic;
  signal Kernel_rematch004_inst_rematch004_in_length         : std_logic_vector(31 downto 0);
  signal Kernel_rematch004_inst_rematch004_in_count          : std_logic_vector(0 downto 0);
  signal Kernel_rematch004_inst_rematch004_in_chars_valid    : std_logic;
  signal Kernel_rematch004_inst_rematch004_in_chars_ready    : std_logic;
  signal Kernel_rematch004_inst_rematch004_in_chars_dvalid   : std_logic;
  signal Kernel_rematch004_inst_rematch004_in_chars_last     : std_logic;
  signal Kernel_rematch004_inst_rematch004_in_chars          : std_logic_vector(31 downto 0);
  signal Kernel_rematch004_inst_rematch004_in_chars_count    : std_logic_vector(2 downto 0);

  signal Kernel_rematch004_inst_rematch004_in_bus_rreq_valid : std_logic;
  signal Kernel_rematch004_inst_rematch004_in_bus_rreq_ready : std_logic;
  signal Kernel_rematch004_inst_rematch004_in_bus_rreq_addr  : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Kernel_rematch004_inst_rematch004_in_bus_rreq_len   : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Kernel_rematch004_inst_rematch004_in_bus_rdat_valid : std_logic;
  signal Kernel_rematch004_inst_rematch004_in_bus_rdat_ready : std_logic;
  signal Kernel_rematch004_inst_rematch004_in_bus_rdat_data  : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Kernel_rematch004_inst_rematch004_in_bus_rdat_last  : std_logic;

  signal Kernel_rematch004_inst_rematch004_in_cmd_valid      : std_logic;
  signal Kernel_rematch004_inst_rematch004_in_cmd_ready      : std_logic;
  signal Kernel_rematch004_inst_rematch004_in_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch004_inst_rematch004_in_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch004_inst_rematch004_in_cmd_ctrl       : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_rematch004_inst_rematch004_in_cmd_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch004_inst_rematch004_in_unl_valid      : std_logic;
  signal Kernel_rematch004_inst_rematch004_in_unl_ready      : std_logic;
  signal Kernel_rematch004_inst_rematch004_in_unl_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch005_inst_rematch005_in_valid          : std_logic;
  signal Kernel_rematch005_inst_rematch005_in_ready          : std_logic;
  signal Kernel_rematch005_inst_rematch005_in_dvalid         : std_logic;
  signal Kernel_rematch005_inst_rematch005_in_last           : std_logic;
  signal Kernel_rematch005_inst_rematch005_in_length         : std_logic_vector(31 downto 0);
  signal Kernel_rematch005_inst_rematch005_in_count          : std_logic_vector(0 downto 0);
  signal Kernel_rematch005_inst_rematch005_in_chars_valid    : std_logic;
  signal Kernel_rematch005_inst_rematch005_in_chars_ready    : std_logic;
  signal Kernel_rematch005_inst_rematch005_in_chars_dvalid   : std_logic;
  signal Kernel_rematch005_inst_rematch005_in_chars_last     : std_logic;
  signal Kernel_rematch005_inst_rematch005_in_chars          : std_logic_vector(31 downto 0);
  signal Kernel_rematch005_inst_rematch005_in_chars_count    : std_logic_vector(2 downto 0);

  signal Kernel_rematch005_inst_rematch005_in_bus_rreq_valid : std_logic;
  signal Kernel_rematch005_inst_rematch005_in_bus_rreq_ready : std_logic;
  signal Kernel_rematch005_inst_rematch005_in_bus_rreq_addr  : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Kernel_rematch005_inst_rematch005_in_bus_rreq_len   : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Kernel_rematch005_inst_rematch005_in_bus_rdat_valid : std_logic;
  signal Kernel_rematch005_inst_rematch005_in_bus_rdat_ready : std_logic;
  signal Kernel_rematch005_inst_rematch005_in_bus_rdat_data  : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Kernel_rematch005_inst_rematch005_in_bus_rdat_last  : std_logic;

  signal Kernel_rematch005_inst_rematch005_in_cmd_valid      : std_logic;
  signal Kernel_rematch005_inst_rematch005_in_cmd_ready      : std_logic;
  signal Kernel_rematch005_inst_rematch005_in_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch005_inst_rematch005_in_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch005_inst_rematch005_in_cmd_ctrl       : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_rematch005_inst_rematch005_in_cmd_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch005_inst_rematch005_in_unl_valid      : std_logic;
  signal Kernel_rematch005_inst_rematch005_in_unl_ready      : std_logic;
  signal Kernel_rematch005_inst_rematch005_in_unl_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch006_inst_rematch006_in_valid          : std_logic;
  signal Kernel_rematch006_inst_rematch006_in_ready          : std_logic;
  signal Kernel_rematch006_inst_rematch006_in_dvalid         : std_logic;
  signal Kernel_rematch006_inst_rematch006_in_last           : std_logic;
  signal Kernel_rematch006_inst_rematch006_in_length         : std_logic_vector(31 downto 0);
  signal Kernel_rematch006_inst_rematch006_in_count          : std_logic_vector(0 downto 0);
  signal Kernel_rematch006_inst_rematch006_in_chars_valid    : std_logic;
  signal Kernel_rematch006_inst_rematch006_in_chars_ready    : std_logic;
  signal Kernel_rematch006_inst_rematch006_in_chars_dvalid   : std_logic;
  signal Kernel_rematch006_inst_rematch006_in_chars_last     : std_logic;
  signal Kernel_rematch006_inst_rematch006_in_chars          : std_logic_vector(31 downto 0);
  signal Kernel_rematch006_inst_rematch006_in_chars_count    : std_logic_vector(2 downto 0);

  signal Kernel_rematch006_inst_rematch006_in_bus_rreq_valid : std_logic;
  signal Kernel_rematch006_inst_rematch006_in_bus_rreq_ready : std_logic;
  signal Kernel_rematch006_inst_rematch006_in_bus_rreq_addr  : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Kernel_rematch006_inst_rematch006_in_bus_rreq_len   : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Kernel_rematch006_inst_rematch006_in_bus_rdat_valid : std_logic;
  signal Kernel_rematch006_inst_rematch006_in_bus_rdat_ready : std_logic;
  signal Kernel_rematch006_inst_rematch006_in_bus_rdat_data  : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Kernel_rematch006_inst_rematch006_in_bus_rdat_last  : std_logic;

  signal Kernel_rematch006_inst_rematch006_in_cmd_valid      : std_logic;
  signal Kernel_rematch006_inst_rematch006_in_cmd_ready      : std_logic;
  signal Kernel_rematch006_inst_rematch006_in_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch006_inst_rematch006_in_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch006_inst_rematch006_in_cmd_ctrl       : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_rematch006_inst_rematch006_in_cmd_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch006_inst_rematch006_in_unl_valid      : std_logic;
  signal Kernel_rematch006_inst_rematch006_in_unl_ready      : std_logic;
  signal Kernel_rematch006_inst_rematch006_in_unl_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch007_inst_rematch007_in_valid          : std_logic;
  signal Kernel_rematch007_inst_rematch007_in_ready          : std_logic;
  signal Kernel_rematch007_inst_rematch007_in_dvalid         : std_logic;
  signal Kernel_rematch007_inst_rematch007_in_last           : std_logic;
  signal Kernel_rematch007_inst_rematch007_in_length         : std_logic_vector(31 downto 0);
  signal Kernel_rematch007_inst_rematch007_in_count          : std_logic_vector(0 downto 0);
  signal Kernel_rematch007_inst_rematch007_in_chars_valid    : std_logic;
  signal Kernel_rematch007_inst_rematch007_in_chars_ready    : std_logic;
  signal Kernel_rematch007_inst_rematch007_in_chars_dvalid   : std_logic;
  signal Kernel_rematch007_inst_rematch007_in_chars_last     : std_logic;
  signal Kernel_rematch007_inst_rematch007_in_chars          : std_logic_vector(31 downto 0);
  signal Kernel_rematch007_inst_rematch007_in_chars_count    : std_logic_vector(2 downto 0);

  signal Kernel_rematch007_inst_rematch007_in_bus_rreq_valid : std_logic;
  signal Kernel_rematch007_inst_rematch007_in_bus_rreq_ready : std_logic;
  signal Kernel_rematch007_inst_rematch007_in_bus_rreq_addr  : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Kernel_rematch007_inst_rematch007_in_bus_rreq_len   : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Kernel_rematch007_inst_rematch007_in_bus_rdat_valid : std_logic;
  signal Kernel_rematch007_inst_rematch007_in_bus_rdat_ready : std_logic;
  signal Kernel_rematch007_inst_rematch007_in_bus_rdat_data  : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Kernel_rematch007_inst_rematch007_in_bus_rdat_last  : std_logic;

  signal Kernel_rematch007_inst_rematch007_in_cmd_valid      : std_logic;
  signal Kernel_rematch007_inst_rematch007_in_cmd_ready      : std_logic;
  signal Kernel_rematch007_inst_rematch007_in_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch007_inst_rematch007_in_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch007_inst_rematch007_in_cmd_ctrl       : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_rematch007_inst_rematch007_in_cmd_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch007_inst_rematch007_in_unl_valid      : std_logic;
  signal Kernel_rematch007_inst_rematch007_in_unl_ready      : std_logic;
  signal Kernel_rematch007_inst_rematch007_in_unl_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch008_inst_rematch008_in_valid          : std_logic;
  signal Kernel_rematch008_inst_rematch008_in_ready          : std_logic;
  signal Kernel_rematch008_inst_rematch008_in_dvalid         : std_logic;
  signal Kernel_rematch008_inst_rematch008_in_last           : std_logic;
  signal Kernel_rematch008_inst_rematch008_in_length         : std_logic_vector(31 downto 0);
  signal Kernel_rematch008_inst_rematch008_in_count          : std_logic_vector(0 downto 0);
  signal Kernel_rematch008_inst_rematch008_in_chars_valid    : std_logic;
  signal Kernel_rematch008_inst_rematch008_in_chars_ready    : std_logic;
  signal Kernel_rematch008_inst_rematch008_in_chars_dvalid   : std_logic;
  signal Kernel_rematch008_inst_rematch008_in_chars_last     : std_logic;
  signal Kernel_rematch008_inst_rematch008_in_chars          : std_logic_vector(31 downto 0);
  signal Kernel_rematch008_inst_rematch008_in_chars_count    : std_logic_vector(2 downto 0);

  signal Kernel_rematch008_inst_rematch008_in_bus_rreq_valid : std_logic;
  signal Kernel_rematch008_inst_rematch008_in_bus_rreq_ready : std_logic;
  signal Kernel_rematch008_inst_rematch008_in_bus_rreq_addr  : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Kernel_rematch008_inst_rematch008_in_bus_rreq_len   : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Kernel_rematch008_inst_rematch008_in_bus_rdat_valid : std_logic;
  signal Kernel_rematch008_inst_rematch008_in_bus_rdat_ready : std_logic;
  signal Kernel_rematch008_inst_rematch008_in_bus_rdat_data  : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Kernel_rematch008_inst_rematch008_in_bus_rdat_last  : std_logic;

  signal Kernel_rematch008_inst_rematch008_in_cmd_valid      : std_logic;
  signal Kernel_rematch008_inst_rematch008_in_cmd_ready      : std_logic;
  signal Kernel_rematch008_inst_rematch008_in_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch008_inst_rematch008_in_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch008_inst_rematch008_in_cmd_ctrl       : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_rematch008_inst_rematch008_in_cmd_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch008_inst_rematch008_in_unl_valid      : std_logic;
  signal Kernel_rematch008_inst_rematch008_in_unl_ready      : std_logic;
  signal Kernel_rematch008_inst_rematch008_in_unl_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch009_inst_rematch009_in_valid          : std_logic;
  signal Kernel_rematch009_inst_rematch009_in_ready          : std_logic;
  signal Kernel_rematch009_inst_rematch009_in_dvalid         : std_logic;
  signal Kernel_rematch009_inst_rematch009_in_last           : std_logic;
  signal Kernel_rematch009_inst_rematch009_in_length         : std_logic_vector(31 downto 0);
  signal Kernel_rematch009_inst_rematch009_in_count          : std_logic_vector(0 downto 0);
  signal Kernel_rematch009_inst_rematch009_in_chars_valid    : std_logic;
  signal Kernel_rematch009_inst_rematch009_in_chars_ready    : std_logic;
  signal Kernel_rematch009_inst_rematch009_in_chars_dvalid   : std_logic;
  signal Kernel_rematch009_inst_rematch009_in_chars_last     : std_logic;
  signal Kernel_rematch009_inst_rematch009_in_chars          : std_logic_vector(31 downto 0);
  signal Kernel_rematch009_inst_rematch009_in_chars_count    : std_logic_vector(2 downto 0);

  signal Kernel_rematch009_inst_rematch009_in_bus_rreq_valid : std_logic;
  signal Kernel_rematch009_inst_rematch009_in_bus_rreq_ready : std_logic;
  signal Kernel_rematch009_inst_rematch009_in_bus_rreq_addr  : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Kernel_rematch009_inst_rematch009_in_bus_rreq_len   : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Kernel_rematch009_inst_rematch009_in_bus_rdat_valid : std_logic;
  signal Kernel_rematch009_inst_rematch009_in_bus_rdat_ready : std_logic;
  signal Kernel_rematch009_inst_rematch009_in_bus_rdat_data  : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Kernel_rematch009_inst_rematch009_in_bus_rdat_last  : std_logic;

  signal Kernel_rematch009_inst_rematch009_in_cmd_valid      : std_logic;
  signal Kernel_rematch009_inst_rematch009_in_cmd_ready      : std_logic;
  signal Kernel_rematch009_inst_rematch009_in_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch009_inst_rematch009_in_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch009_inst_rematch009_in_cmd_ctrl       : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_rematch009_inst_rematch009_in_cmd_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch009_inst_rematch009_in_unl_valid      : std_logic;
  signal Kernel_rematch009_inst_rematch009_in_unl_ready      : std_logic;
  signal Kernel_rematch009_inst_rematch009_in_unl_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch010_inst_rematch010_in_valid          : std_logic;
  signal Kernel_rematch010_inst_rematch010_in_ready          : std_logic;
  signal Kernel_rematch010_inst_rematch010_in_dvalid         : std_logic;
  signal Kernel_rematch010_inst_rematch010_in_last           : std_logic;
  signal Kernel_rematch010_inst_rematch010_in_length         : std_logic_vector(31 downto 0);
  signal Kernel_rematch010_inst_rematch010_in_count          : std_logic_vector(0 downto 0);
  signal Kernel_rematch010_inst_rematch010_in_chars_valid    : std_logic;
  signal Kernel_rematch010_inst_rematch010_in_chars_ready    : std_logic;
  signal Kernel_rematch010_inst_rematch010_in_chars_dvalid   : std_logic;
  signal Kernel_rematch010_inst_rematch010_in_chars_last     : std_logic;
  signal Kernel_rematch010_inst_rematch010_in_chars          : std_logic_vector(31 downto 0);
  signal Kernel_rematch010_inst_rematch010_in_chars_count    : std_logic_vector(2 downto 0);

  signal Kernel_rematch010_inst_rematch010_in_bus_rreq_valid : std_logic;
  signal Kernel_rematch010_inst_rematch010_in_bus_rreq_ready : std_logic;
  signal Kernel_rematch010_inst_rematch010_in_bus_rreq_addr  : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Kernel_rematch010_inst_rematch010_in_bus_rreq_len   : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Kernel_rematch010_inst_rematch010_in_bus_rdat_valid : std_logic;
  signal Kernel_rematch010_inst_rematch010_in_bus_rdat_ready : std_logic;
  signal Kernel_rematch010_inst_rematch010_in_bus_rdat_data  : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Kernel_rematch010_inst_rematch010_in_bus_rdat_last  : std_logic;

  signal Kernel_rematch010_inst_rematch010_in_cmd_valid      : std_logic;
  signal Kernel_rematch010_inst_rematch010_in_cmd_ready      : std_logic;
  signal Kernel_rematch010_inst_rematch010_in_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch010_inst_rematch010_in_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch010_inst_rematch010_in_cmd_ctrl       : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_rematch010_inst_rematch010_in_cmd_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch010_inst_rematch010_in_unl_valid      : std_logic;
  signal Kernel_rematch010_inst_rematch010_in_unl_ready      : std_logic;
  signal Kernel_rematch010_inst_rematch010_in_unl_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch011_inst_rematch011_in_valid          : std_logic;
  signal Kernel_rematch011_inst_rematch011_in_ready          : std_logic;
  signal Kernel_rematch011_inst_rematch011_in_dvalid         : std_logic;
  signal Kernel_rematch011_inst_rematch011_in_last           : std_logic;
  signal Kernel_rematch011_inst_rematch011_in_length         : std_logic_vector(31 downto 0);
  signal Kernel_rematch011_inst_rematch011_in_count          : std_logic_vector(0 downto 0);
  signal Kernel_rematch011_inst_rematch011_in_chars_valid    : std_logic;
  signal Kernel_rematch011_inst_rematch011_in_chars_ready    : std_logic;
  signal Kernel_rematch011_inst_rematch011_in_chars_dvalid   : std_logic;
  signal Kernel_rematch011_inst_rematch011_in_chars_last     : std_logic;
  signal Kernel_rematch011_inst_rematch011_in_chars          : std_logic_vector(31 downto 0);
  signal Kernel_rematch011_inst_rematch011_in_chars_count    : std_logic_vector(2 downto 0);

  signal Kernel_rematch011_inst_rematch011_in_bus_rreq_valid : std_logic;
  signal Kernel_rematch011_inst_rematch011_in_bus_rreq_ready : std_logic;
  signal Kernel_rematch011_inst_rematch011_in_bus_rreq_addr  : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Kernel_rematch011_inst_rematch011_in_bus_rreq_len   : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Kernel_rematch011_inst_rematch011_in_bus_rdat_valid : std_logic;
  signal Kernel_rematch011_inst_rematch011_in_bus_rdat_ready : std_logic;
  signal Kernel_rematch011_inst_rematch011_in_bus_rdat_data  : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Kernel_rematch011_inst_rematch011_in_bus_rdat_last  : std_logic;

  signal Kernel_rematch011_inst_rematch011_in_cmd_valid      : std_logic;
  signal Kernel_rematch011_inst_rematch011_in_cmd_ready      : std_logic;
  signal Kernel_rematch011_inst_rematch011_in_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch011_inst_rematch011_in_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch011_inst_rematch011_in_cmd_ctrl       : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_rematch011_inst_rematch011_in_cmd_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch011_inst_rematch011_in_unl_valid      : std_logic;
  signal Kernel_rematch011_inst_rematch011_in_unl_ready      : std_logic;
  signal Kernel_rematch011_inst_rematch011_in_unl_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch012_inst_rematch012_in_valid          : std_logic;
  signal Kernel_rematch012_inst_rematch012_in_ready          : std_logic;
  signal Kernel_rematch012_inst_rematch012_in_dvalid         : std_logic;
  signal Kernel_rematch012_inst_rematch012_in_last           : std_logic;
  signal Kernel_rematch012_inst_rematch012_in_length         : std_logic_vector(31 downto 0);
  signal Kernel_rematch012_inst_rematch012_in_count          : std_logic_vector(0 downto 0);
  signal Kernel_rematch012_inst_rematch012_in_chars_valid    : std_logic;
  signal Kernel_rematch012_inst_rematch012_in_chars_ready    : std_logic;
  signal Kernel_rematch012_inst_rematch012_in_chars_dvalid   : std_logic;
  signal Kernel_rematch012_inst_rematch012_in_chars_last     : std_logic;
  signal Kernel_rematch012_inst_rematch012_in_chars          : std_logic_vector(31 downto 0);
  signal Kernel_rematch012_inst_rematch012_in_chars_count    : std_logic_vector(2 downto 0);

  signal Kernel_rematch012_inst_rematch012_in_bus_rreq_valid : std_logic;
  signal Kernel_rematch012_inst_rematch012_in_bus_rreq_ready : std_logic;
  signal Kernel_rematch012_inst_rematch012_in_bus_rreq_addr  : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Kernel_rematch012_inst_rematch012_in_bus_rreq_len   : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Kernel_rematch012_inst_rematch012_in_bus_rdat_valid : std_logic;
  signal Kernel_rematch012_inst_rematch012_in_bus_rdat_ready : std_logic;
  signal Kernel_rematch012_inst_rematch012_in_bus_rdat_data  : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Kernel_rematch012_inst_rematch012_in_bus_rdat_last  : std_logic;

  signal Kernel_rematch012_inst_rematch012_in_cmd_valid      : std_logic;
  signal Kernel_rematch012_inst_rematch012_in_cmd_ready      : std_logic;
  signal Kernel_rematch012_inst_rematch012_in_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch012_inst_rematch012_in_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch012_inst_rematch012_in_cmd_ctrl       : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_rematch012_inst_rematch012_in_cmd_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch012_inst_rematch012_in_unl_valid      : std_logic;
  signal Kernel_rematch012_inst_rematch012_in_unl_ready      : std_logic;
  signal Kernel_rematch012_inst_rematch012_in_unl_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch013_inst_rematch013_in_valid          : std_logic;
  signal Kernel_rematch013_inst_rematch013_in_ready          : std_logic;
  signal Kernel_rematch013_inst_rematch013_in_dvalid         : std_logic;
  signal Kernel_rematch013_inst_rematch013_in_last           : std_logic;
  signal Kernel_rematch013_inst_rematch013_in_length         : std_logic_vector(31 downto 0);
  signal Kernel_rematch013_inst_rematch013_in_count          : std_logic_vector(0 downto 0);
  signal Kernel_rematch013_inst_rematch013_in_chars_valid    : std_logic;
  signal Kernel_rematch013_inst_rematch013_in_chars_ready    : std_logic;
  signal Kernel_rematch013_inst_rematch013_in_chars_dvalid   : std_logic;
  signal Kernel_rematch013_inst_rematch013_in_chars_last     : std_logic;
  signal Kernel_rematch013_inst_rematch013_in_chars          : std_logic_vector(31 downto 0);
  signal Kernel_rematch013_inst_rematch013_in_chars_count    : std_logic_vector(2 downto 0);

  signal Kernel_rematch013_inst_rematch013_in_bus_rreq_valid : std_logic;
  signal Kernel_rematch013_inst_rematch013_in_bus_rreq_ready : std_logic;
  signal Kernel_rematch013_inst_rematch013_in_bus_rreq_addr  : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Kernel_rematch013_inst_rematch013_in_bus_rreq_len   : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Kernel_rematch013_inst_rematch013_in_bus_rdat_valid : std_logic;
  signal Kernel_rematch013_inst_rematch013_in_bus_rdat_ready : std_logic;
  signal Kernel_rematch013_inst_rematch013_in_bus_rdat_data  : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Kernel_rematch013_inst_rematch013_in_bus_rdat_last  : std_logic;

  signal Kernel_rematch013_inst_rematch013_in_cmd_valid      : std_logic;
  signal Kernel_rematch013_inst_rematch013_in_cmd_ready      : std_logic;
  signal Kernel_rematch013_inst_rematch013_in_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch013_inst_rematch013_in_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch013_inst_rematch013_in_cmd_ctrl       : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_rematch013_inst_rematch013_in_cmd_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch013_inst_rematch013_in_unl_valid      : std_logic;
  signal Kernel_rematch013_inst_rematch013_in_unl_ready      : std_logic;
  signal Kernel_rematch013_inst_rematch013_in_unl_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch014_inst_rematch014_in_valid          : std_logic;
  signal Kernel_rematch014_inst_rematch014_in_ready          : std_logic;
  signal Kernel_rematch014_inst_rematch014_in_dvalid         : std_logic;
  signal Kernel_rematch014_inst_rematch014_in_last           : std_logic;
  signal Kernel_rematch014_inst_rematch014_in_length         : std_logic_vector(31 downto 0);
  signal Kernel_rematch014_inst_rematch014_in_count          : std_logic_vector(0 downto 0);
  signal Kernel_rematch014_inst_rematch014_in_chars_valid    : std_logic;
  signal Kernel_rematch014_inst_rematch014_in_chars_ready    : std_logic;
  signal Kernel_rematch014_inst_rematch014_in_chars_dvalid   : std_logic;
  signal Kernel_rematch014_inst_rematch014_in_chars_last     : std_logic;
  signal Kernel_rematch014_inst_rematch014_in_chars          : std_logic_vector(31 downto 0);
  signal Kernel_rematch014_inst_rematch014_in_chars_count    : std_logic_vector(2 downto 0);

  signal Kernel_rematch014_inst_rematch014_in_bus_rreq_valid : std_logic;
  signal Kernel_rematch014_inst_rematch014_in_bus_rreq_ready : std_logic;
  signal Kernel_rematch014_inst_rematch014_in_bus_rreq_addr  : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Kernel_rematch014_inst_rematch014_in_bus_rreq_len   : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Kernel_rematch014_inst_rematch014_in_bus_rdat_valid : std_logic;
  signal Kernel_rematch014_inst_rematch014_in_bus_rdat_ready : std_logic;
  signal Kernel_rematch014_inst_rematch014_in_bus_rdat_data  : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Kernel_rematch014_inst_rematch014_in_bus_rdat_last  : std_logic;

  signal Kernel_rematch014_inst_rematch014_in_cmd_valid      : std_logic;
  signal Kernel_rematch014_inst_rematch014_in_cmd_ready      : std_logic;
  signal Kernel_rematch014_inst_rematch014_in_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch014_inst_rematch014_in_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch014_inst_rematch014_in_cmd_ctrl       : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_rematch014_inst_rematch014_in_cmd_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch014_inst_rematch014_in_unl_valid      : std_logic;
  signal Kernel_rematch014_inst_rematch014_in_unl_ready      : std_logic;
  signal Kernel_rematch014_inst_rematch014_in_unl_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch015_inst_rematch015_in_valid          : std_logic;
  signal Kernel_rematch015_inst_rematch015_in_ready          : std_logic;
  signal Kernel_rematch015_inst_rematch015_in_dvalid         : std_logic;
  signal Kernel_rematch015_inst_rematch015_in_last           : std_logic;
  signal Kernel_rematch015_inst_rematch015_in_length         : std_logic_vector(31 downto 0);
  signal Kernel_rematch015_inst_rematch015_in_count          : std_logic_vector(0 downto 0);
  signal Kernel_rematch015_inst_rematch015_in_chars_valid    : std_logic;
  signal Kernel_rematch015_inst_rematch015_in_chars_ready    : std_logic;
  signal Kernel_rematch015_inst_rematch015_in_chars_dvalid   : std_logic;
  signal Kernel_rematch015_inst_rematch015_in_chars_last     : std_logic;
  signal Kernel_rematch015_inst_rematch015_in_chars          : std_logic_vector(31 downto 0);
  signal Kernel_rematch015_inst_rematch015_in_chars_count    : std_logic_vector(2 downto 0);

  signal Kernel_rematch015_inst_rematch015_in_bus_rreq_valid : std_logic;
  signal Kernel_rematch015_inst_rematch015_in_bus_rreq_ready : std_logic;
  signal Kernel_rematch015_inst_rematch015_in_bus_rreq_addr  : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Kernel_rematch015_inst_rematch015_in_bus_rreq_len   : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Kernel_rematch015_inst_rematch015_in_bus_rdat_valid : std_logic;
  signal Kernel_rematch015_inst_rematch015_in_bus_rdat_ready : std_logic;
  signal Kernel_rematch015_inst_rematch015_in_bus_rdat_data  : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Kernel_rematch015_inst_rematch015_in_bus_rdat_last  : std_logic;

  signal Kernel_rematch015_inst_rematch015_in_cmd_valid      : std_logic;
  signal Kernel_rematch015_inst_rematch015_in_cmd_ready      : std_logic;
  signal Kernel_rematch015_inst_rematch015_in_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch015_inst_rematch015_in_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Kernel_rematch015_inst_rematch015_in_cmd_ctrl       : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal Kernel_rematch015_inst_rematch015_in_cmd_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Kernel_rematch015_inst_rematch015_in_unl_valid      : std_logic;
  signal Kernel_rematch015_inst_rematch015_in_unl_ready      : std_logic;
  signal Kernel_rematch015_inst_rematch015_in_unl_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_valid           : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_ready           : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_addr            : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_len             : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_valid           : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_ready           : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_data            : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_last            : std_logic;

  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid : std_logic_vector(15 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready : std_logic_vector(15 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr  : std_logic_vector(16*BUS_ADDR_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len   : std_logic_vector(16*BUS_LEN_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid : std_logic_vector(15 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready : std_logic_vector(15 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data  : std_logic_vector(16*BUS_DATA_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last  : std_logic_vector(15 downto 0);

begin
  Kernel_Nucleus_inst : Kernel_Nucleus
    generic map (
      INDEX_WIDTH                  => INDEX_WIDTH,
      TAG_WIDTH                    => TAG_WIDTH,
      REMATCH000_IN_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
      REMATCH001_IN_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
      REMATCH002_IN_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
      REMATCH003_IN_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
      REMATCH004_IN_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
      REMATCH005_IN_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
      REMATCH006_IN_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
      REMATCH007_IN_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
      REMATCH008_IN_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
      REMATCH009_IN_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
      REMATCH010_IN_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
      REMATCH011_IN_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
      REMATCH012_IN_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
      REMATCH013_IN_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
      REMATCH014_IN_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
      REMATCH015_IN_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH
    )
    port map (
      kcd_clk                    => kcd_clk,
      kcd_reset                  => kcd_reset,
      mmio_awvalid               => Kernel_Nucleus_inst_mmio_awvalid,
      mmio_awready               => Kernel_Nucleus_inst_mmio_awready,
      mmio_awaddr                => Kernel_Nucleus_inst_mmio_awaddr,
      mmio_wvalid                => Kernel_Nucleus_inst_mmio_wvalid,
      mmio_wready                => Kernel_Nucleus_inst_mmio_wready,
      mmio_wdata                 => Kernel_Nucleus_inst_mmio_wdata,
      mmio_wstrb                 => Kernel_Nucleus_inst_mmio_wstrb,
      mmio_bvalid                => Kernel_Nucleus_inst_mmio_bvalid,
      mmio_bready                => Kernel_Nucleus_inst_mmio_bready,
      mmio_bresp                 => Kernel_Nucleus_inst_mmio_bresp,
      mmio_arvalid               => Kernel_Nucleus_inst_mmio_arvalid,
      mmio_arready               => Kernel_Nucleus_inst_mmio_arready,
      mmio_araddr                => Kernel_Nucleus_inst_mmio_araddr,
      mmio_rvalid                => Kernel_Nucleus_inst_mmio_rvalid,
      mmio_rready                => Kernel_Nucleus_inst_mmio_rready,
      mmio_rdata                 => Kernel_Nucleus_inst_mmio_rdata,
      mmio_rresp                 => Kernel_Nucleus_inst_mmio_rresp,
      rematch000_in_valid        => Kernel_Nucleus_inst_rematch000_in_valid,
      rematch000_in_ready        => Kernel_Nucleus_inst_rematch000_in_ready,
      rematch000_in_dvalid       => Kernel_Nucleus_inst_rematch000_in_dvalid,
      rematch000_in_last         => Kernel_Nucleus_inst_rematch000_in_last,
      rematch000_in_length       => Kernel_Nucleus_inst_rematch000_in_length,
      rematch000_in_count        => Kernel_Nucleus_inst_rematch000_in_count,
      rematch000_in_chars_valid  => Kernel_Nucleus_inst_rematch000_in_chars_valid,
      rematch000_in_chars_ready  => Kernel_Nucleus_inst_rematch000_in_chars_ready,
      rematch000_in_chars_dvalid => Kernel_Nucleus_inst_rematch000_in_chars_dvalid,
      rematch000_in_chars_last   => Kernel_Nucleus_inst_rematch000_in_chars_last,
      rematch000_in_chars        => Kernel_Nucleus_inst_rematch000_in_chars,
      rematch000_in_chars_count  => Kernel_Nucleus_inst_rematch000_in_chars_count,
      rematch000_in_unl_valid    => Kernel_Nucleus_inst_rematch000_in_unl_valid,
      rematch000_in_unl_ready    => Kernel_Nucleus_inst_rematch000_in_unl_ready,
      rematch000_in_unl_tag      => Kernel_Nucleus_inst_rematch000_in_unl_tag,
      rematch000_in_cmd_valid    => Kernel_Nucleus_inst_rematch000_in_cmd_valid,
      rematch000_in_cmd_ready    => Kernel_Nucleus_inst_rematch000_in_cmd_ready,
      rematch000_in_cmd_firstIdx => Kernel_Nucleus_inst_rematch000_in_cmd_firstIdx,
      rematch000_in_cmd_lastIdx  => Kernel_Nucleus_inst_rematch000_in_cmd_lastIdx,
      rematch000_in_cmd_ctrl     => Kernel_Nucleus_inst_rematch000_in_cmd_ctrl,
      rematch000_in_cmd_tag      => Kernel_Nucleus_inst_rematch000_in_cmd_tag,
      rematch001_in_valid        => Kernel_Nucleus_inst_rematch001_in_valid,
      rematch001_in_ready        => Kernel_Nucleus_inst_rematch001_in_ready,
      rematch001_in_dvalid       => Kernel_Nucleus_inst_rematch001_in_dvalid,
      rematch001_in_last         => Kernel_Nucleus_inst_rematch001_in_last,
      rematch001_in_length       => Kernel_Nucleus_inst_rematch001_in_length,
      rematch001_in_count        => Kernel_Nucleus_inst_rematch001_in_count,
      rematch001_in_chars_valid  => Kernel_Nucleus_inst_rematch001_in_chars_valid,
      rematch001_in_chars_ready  => Kernel_Nucleus_inst_rematch001_in_chars_ready,
      rematch001_in_chars_dvalid => Kernel_Nucleus_inst_rematch001_in_chars_dvalid,
      rematch001_in_chars_last   => Kernel_Nucleus_inst_rematch001_in_chars_last,
      rematch001_in_chars        => Kernel_Nucleus_inst_rematch001_in_chars,
      rematch001_in_chars_count  => Kernel_Nucleus_inst_rematch001_in_chars_count,
      rematch001_in_unl_valid    => Kernel_Nucleus_inst_rematch001_in_unl_valid,
      rematch001_in_unl_ready    => Kernel_Nucleus_inst_rematch001_in_unl_ready,
      rematch001_in_unl_tag      => Kernel_Nucleus_inst_rematch001_in_unl_tag,
      rematch001_in_cmd_valid    => Kernel_Nucleus_inst_rematch001_in_cmd_valid,
      rematch001_in_cmd_ready    => Kernel_Nucleus_inst_rematch001_in_cmd_ready,
      rematch001_in_cmd_firstIdx => Kernel_Nucleus_inst_rematch001_in_cmd_firstIdx,
      rematch001_in_cmd_lastIdx  => Kernel_Nucleus_inst_rematch001_in_cmd_lastIdx,
      rematch001_in_cmd_ctrl     => Kernel_Nucleus_inst_rematch001_in_cmd_ctrl,
      rematch001_in_cmd_tag      => Kernel_Nucleus_inst_rematch001_in_cmd_tag,
      rematch002_in_valid        => Kernel_Nucleus_inst_rematch002_in_valid,
      rematch002_in_ready        => Kernel_Nucleus_inst_rematch002_in_ready,
      rematch002_in_dvalid       => Kernel_Nucleus_inst_rematch002_in_dvalid,
      rematch002_in_last         => Kernel_Nucleus_inst_rematch002_in_last,
      rematch002_in_length       => Kernel_Nucleus_inst_rematch002_in_length,
      rematch002_in_count        => Kernel_Nucleus_inst_rematch002_in_count,
      rematch002_in_chars_valid  => Kernel_Nucleus_inst_rematch002_in_chars_valid,
      rematch002_in_chars_ready  => Kernel_Nucleus_inst_rematch002_in_chars_ready,
      rematch002_in_chars_dvalid => Kernel_Nucleus_inst_rematch002_in_chars_dvalid,
      rematch002_in_chars_last   => Kernel_Nucleus_inst_rematch002_in_chars_last,
      rematch002_in_chars        => Kernel_Nucleus_inst_rematch002_in_chars,
      rematch002_in_chars_count  => Kernel_Nucleus_inst_rematch002_in_chars_count,
      rematch002_in_unl_valid    => Kernel_Nucleus_inst_rematch002_in_unl_valid,
      rematch002_in_unl_ready    => Kernel_Nucleus_inst_rematch002_in_unl_ready,
      rematch002_in_unl_tag      => Kernel_Nucleus_inst_rematch002_in_unl_tag,
      rematch002_in_cmd_valid    => Kernel_Nucleus_inst_rematch002_in_cmd_valid,
      rematch002_in_cmd_ready    => Kernel_Nucleus_inst_rematch002_in_cmd_ready,
      rematch002_in_cmd_firstIdx => Kernel_Nucleus_inst_rematch002_in_cmd_firstIdx,
      rematch002_in_cmd_lastIdx  => Kernel_Nucleus_inst_rematch002_in_cmd_lastIdx,
      rematch002_in_cmd_ctrl     => Kernel_Nucleus_inst_rematch002_in_cmd_ctrl,
      rematch002_in_cmd_tag      => Kernel_Nucleus_inst_rematch002_in_cmd_tag,
      rematch003_in_valid        => Kernel_Nucleus_inst_rematch003_in_valid,
      rematch003_in_ready        => Kernel_Nucleus_inst_rematch003_in_ready,
      rematch003_in_dvalid       => Kernel_Nucleus_inst_rematch003_in_dvalid,
      rematch003_in_last         => Kernel_Nucleus_inst_rematch003_in_last,
      rematch003_in_length       => Kernel_Nucleus_inst_rematch003_in_length,
      rematch003_in_count        => Kernel_Nucleus_inst_rematch003_in_count,
      rematch003_in_chars_valid  => Kernel_Nucleus_inst_rematch003_in_chars_valid,
      rematch003_in_chars_ready  => Kernel_Nucleus_inst_rematch003_in_chars_ready,
      rematch003_in_chars_dvalid => Kernel_Nucleus_inst_rematch003_in_chars_dvalid,
      rematch003_in_chars_last   => Kernel_Nucleus_inst_rematch003_in_chars_last,
      rematch003_in_chars        => Kernel_Nucleus_inst_rematch003_in_chars,
      rematch003_in_chars_count  => Kernel_Nucleus_inst_rematch003_in_chars_count,
      rematch003_in_unl_valid    => Kernel_Nucleus_inst_rematch003_in_unl_valid,
      rematch003_in_unl_ready    => Kernel_Nucleus_inst_rematch003_in_unl_ready,
      rematch003_in_unl_tag      => Kernel_Nucleus_inst_rematch003_in_unl_tag,
      rematch003_in_cmd_valid    => Kernel_Nucleus_inst_rematch003_in_cmd_valid,
      rematch003_in_cmd_ready    => Kernel_Nucleus_inst_rematch003_in_cmd_ready,
      rematch003_in_cmd_firstIdx => Kernel_Nucleus_inst_rematch003_in_cmd_firstIdx,
      rematch003_in_cmd_lastIdx  => Kernel_Nucleus_inst_rematch003_in_cmd_lastIdx,
      rematch003_in_cmd_ctrl     => Kernel_Nucleus_inst_rematch003_in_cmd_ctrl,
      rematch003_in_cmd_tag      => Kernel_Nucleus_inst_rematch003_in_cmd_tag,
      rematch004_in_valid        => Kernel_Nucleus_inst_rematch004_in_valid,
      rematch004_in_ready        => Kernel_Nucleus_inst_rematch004_in_ready,
      rematch004_in_dvalid       => Kernel_Nucleus_inst_rematch004_in_dvalid,
      rematch004_in_last         => Kernel_Nucleus_inst_rematch004_in_last,
      rematch004_in_length       => Kernel_Nucleus_inst_rematch004_in_length,
      rematch004_in_count        => Kernel_Nucleus_inst_rematch004_in_count,
      rematch004_in_chars_valid  => Kernel_Nucleus_inst_rematch004_in_chars_valid,
      rematch004_in_chars_ready  => Kernel_Nucleus_inst_rematch004_in_chars_ready,
      rematch004_in_chars_dvalid => Kernel_Nucleus_inst_rematch004_in_chars_dvalid,
      rematch004_in_chars_last   => Kernel_Nucleus_inst_rematch004_in_chars_last,
      rematch004_in_chars        => Kernel_Nucleus_inst_rematch004_in_chars,
      rematch004_in_chars_count  => Kernel_Nucleus_inst_rematch004_in_chars_count,
      rematch004_in_unl_valid    => Kernel_Nucleus_inst_rematch004_in_unl_valid,
      rematch004_in_unl_ready    => Kernel_Nucleus_inst_rematch004_in_unl_ready,
      rematch004_in_unl_tag      => Kernel_Nucleus_inst_rematch004_in_unl_tag,
      rematch004_in_cmd_valid    => Kernel_Nucleus_inst_rematch004_in_cmd_valid,
      rematch004_in_cmd_ready    => Kernel_Nucleus_inst_rematch004_in_cmd_ready,
      rematch004_in_cmd_firstIdx => Kernel_Nucleus_inst_rematch004_in_cmd_firstIdx,
      rematch004_in_cmd_lastIdx  => Kernel_Nucleus_inst_rematch004_in_cmd_lastIdx,
      rematch004_in_cmd_ctrl     => Kernel_Nucleus_inst_rematch004_in_cmd_ctrl,
      rematch004_in_cmd_tag      => Kernel_Nucleus_inst_rematch004_in_cmd_tag,
      rematch005_in_valid        => Kernel_Nucleus_inst_rematch005_in_valid,
      rematch005_in_ready        => Kernel_Nucleus_inst_rematch005_in_ready,
      rematch005_in_dvalid       => Kernel_Nucleus_inst_rematch005_in_dvalid,
      rematch005_in_last         => Kernel_Nucleus_inst_rematch005_in_last,
      rematch005_in_length       => Kernel_Nucleus_inst_rematch005_in_length,
      rematch005_in_count        => Kernel_Nucleus_inst_rematch005_in_count,
      rematch005_in_chars_valid  => Kernel_Nucleus_inst_rematch005_in_chars_valid,
      rematch005_in_chars_ready  => Kernel_Nucleus_inst_rematch005_in_chars_ready,
      rematch005_in_chars_dvalid => Kernel_Nucleus_inst_rematch005_in_chars_dvalid,
      rematch005_in_chars_last   => Kernel_Nucleus_inst_rematch005_in_chars_last,
      rematch005_in_chars        => Kernel_Nucleus_inst_rematch005_in_chars,
      rematch005_in_chars_count  => Kernel_Nucleus_inst_rematch005_in_chars_count,
      rematch005_in_unl_valid    => Kernel_Nucleus_inst_rematch005_in_unl_valid,
      rematch005_in_unl_ready    => Kernel_Nucleus_inst_rematch005_in_unl_ready,
      rematch005_in_unl_tag      => Kernel_Nucleus_inst_rematch005_in_unl_tag,
      rematch005_in_cmd_valid    => Kernel_Nucleus_inst_rematch005_in_cmd_valid,
      rematch005_in_cmd_ready    => Kernel_Nucleus_inst_rematch005_in_cmd_ready,
      rematch005_in_cmd_firstIdx => Kernel_Nucleus_inst_rematch005_in_cmd_firstIdx,
      rematch005_in_cmd_lastIdx  => Kernel_Nucleus_inst_rematch005_in_cmd_lastIdx,
      rematch005_in_cmd_ctrl     => Kernel_Nucleus_inst_rematch005_in_cmd_ctrl,
      rematch005_in_cmd_tag      => Kernel_Nucleus_inst_rematch005_in_cmd_tag,
      rematch006_in_valid        => Kernel_Nucleus_inst_rematch006_in_valid,
      rematch006_in_ready        => Kernel_Nucleus_inst_rematch006_in_ready,
      rematch006_in_dvalid       => Kernel_Nucleus_inst_rematch006_in_dvalid,
      rematch006_in_last         => Kernel_Nucleus_inst_rematch006_in_last,
      rematch006_in_length       => Kernel_Nucleus_inst_rematch006_in_length,
      rematch006_in_count        => Kernel_Nucleus_inst_rematch006_in_count,
      rematch006_in_chars_valid  => Kernel_Nucleus_inst_rematch006_in_chars_valid,
      rematch006_in_chars_ready  => Kernel_Nucleus_inst_rematch006_in_chars_ready,
      rematch006_in_chars_dvalid => Kernel_Nucleus_inst_rematch006_in_chars_dvalid,
      rematch006_in_chars_last   => Kernel_Nucleus_inst_rematch006_in_chars_last,
      rematch006_in_chars        => Kernel_Nucleus_inst_rematch006_in_chars,
      rematch006_in_chars_count  => Kernel_Nucleus_inst_rematch006_in_chars_count,
      rematch006_in_unl_valid    => Kernel_Nucleus_inst_rematch006_in_unl_valid,
      rematch006_in_unl_ready    => Kernel_Nucleus_inst_rematch006_in_unl_ready,
      rematch006_in_unl_tag      => Kernel_Nucleus_inst_rematch006_in_unl_tag,
      rematch006_in_cmd_valid    => Kernel_Nucleus_inst_rematch006_in_cmd_valid,
      rematch006_in_cmd_ready    => Kernel_Nucleus_inst_rematch006_in_cmd_ready,
      rematch006_in_cmd_firstIdx => Kernel_Nucleus_inst_rematch006_in_cmd_firstIdx,
      rematch006_in_cmd_lastIdx  => Kernel_Nucleus_inst_rematch006_in_cmd_lastIdx,
      rematch006_in_cmd_ctrl     => Kernel_Nucleus_inst_rematch006_in_cmd_ctrl,
      rematch006_in_cmd_tag      => Kernel_Nucleus_inst_rematch006_in_cmd_tag,
      rematch007_in_valid        => Kernel_Nucleus_inst_rematch007_in_valid,
      rematch007_in_ready        => Kernel_Nucleus_inst_rematch007_in_ready,
      rematch007_in_dvalid       => Kernel_Nucleus_inst_rematch007_in_dvalid,
      rematch007_in_last         => Kernel_Nucleus_inst_rematch007_in_last,
      rematch007_in_length       => Kernel_Nucleus_inst_rematch007_in_length,
      rematch007_in_count        => Kernel_Nucleus_inst_rematch007_in_count,
      rematch007_in_chars_valid  => Kernel_Nucleus_inst_rematch007_in_chars_valid,
      rematch007_in_chars_ready  => Kernel_Nucleus_inst_rematch007_in_chars_ready,
      rematch007_in_chars_dvalid => Kernel_Nucleus_inst_rematch007_in_chars_dvalid,
      rematch007_in_chars_last   => Kernel_Nucleus_inst_rematch007_in_chars_last,
      rematch007_in_chars        => Kernel_Nucleus_inst_rematch007_in_chars,
      rematch007_in_chars_count  => Kernel_Nucleus_inst_rematch007_in_chars_count,
      rematch007_in_unl_valid    => Kernel_Nucleus_inst_rematch007_in_unl_valid,
      rematch007_in_unl_ready    => Kernel_Nucleus_inst_rematch007_in_unl_ready,
      rematch007_in_unl_tag      => Kernel_Nucleus_inst_rematch007_in_unl_tag,
      rematch007_in_cmd_valid    => Kernel_Nucleus_inst_rematch007_in_cmd_valid,
      rematch007_in_cmd_ready    => Kernel_Nucleus_inst_rematch007_in_cmd_ready,
      rematch007_in_cmd_firstIdx => Kernel_Nucleus_inst_rematch007_in_cmd_firstIdx,
      rematch007_in_cmd_lastIdx  => Kernel_Nucleus_inst_rematch007_in_cmd_lastIdx,
      rematch007_in_cmd_ctrl     => Kernel_Nucleus_inst_rematch007_in_cmd_ctrl,
      rematch007_in_cmd_tag      => Kernel_Nucleus_inst_rematch007_in_cmd_tag,
      rematch008_in_valid        => Kernel_Nucleus_inst_rematch008_in_valid,
      rematch008_in_ready        => Kernel_Nucleus_inst_rematch008_in_ready,
      rematch008_in_dvalid       => Kernel_Nucleus_inst_rematch008_in_dvalid,
      rematch008_in_last         => Kernel_Nucleus_inst_rematch008_in_last,
      rematch008_in_length       => Kernel_Nucleus_inst_rematch008_in_length,
      rematch008_in_count        => Kernel_Nucleus_inst_rematch008_in_count,
      rematch008_in_chars_valid  => Kernel_Nucleus_inst_rematch008_in_chars_valid,
      rematch008_in_chars_ready  => Kernel_Nucleus_inst_rematch008_in_chars_ready,
      rematch008_in_chars_dvalid => Kernel_Nucleus_inst_rematch008_in_chars_dvalid,
      rematch008_in_chars_last   => Kernel_Nucleus_inst_rematch008_in_chars_last,
      rematch008_in_chars        => Kernel_Nucleus_inst_rematch008_in_chars,
      rematch008_in_chars_count  => Kernel_Nucleus_inst_rematch008_in_chars_count,
      rematch008_in_unl_valid    => Kernel_Nucleus_inst_rematch008_in_unl_valid,
      rematch008_in_unl_ready    => Kernel_Nucleus_inst_rematch008_in_unl_ready,
      rematch008_in_unl_tag      => Kernel_Nucleus_inst_rematch008_in_unl_tag,
      rematch008_in_cmd_valid    => Kernel_Nucleus_inst_rematch008_in_cmd_valid,
      rematch008_in_cmd_ready    => Kernel_Nucleus_inst_rematch008_in_cmd_ready,
      rematch008_in_cmd_firstIdx => Kernel_Nucleus_inst_rematch008_in_cmd_firstIdx,
      rematch008_in_cmd_lastIdx  => Kernel_Nucleus_inst_rematch008_in_cmd_lastIdx,
      rematch008_in_cmd_ctrl     => Kernel_Nucleus_inst_rematch008_in_cmd_ctrl,
      rematch008_in_cmd_tag      => Kernel_Nucleus_inst_rematch008_in_cmd_tag,
      rematch009_in_valid        => Kernel_Nucleus_inst_rematch009_in_valid,
      rematch009_in_ready        => Kernel_Nucleus_inst_rematch009_in_ready,
      rematch009_in_dvalid       => Kernel_Nucleus_inst_rematch009_in_dvalid,
      rematch009_in_last         => Kernel_Nucleus_inst_rematch009_in_last,
      rematch009_in_length       => Kernel_Nucleus_inst_rematch009_in_length,
      rematch009_in_count        => Kernel_Nucleus_inst_rematch009_in_count,
      rematch009_in_chars_valid  => Kernel_Nucleus_inst_rematch009_in_chars_valid,
      rematch009_in_chars_ready  => Kernel_Nucleus_inst_rematch009_in_chars_ready,
      rematch009_in_chars_dvalid => Kernel_Nucleus_inst_rematch009_in_chars_dvalid,
      rematch009_in_chars_last   => Kernel_Nucleus_inst_rematch009_in_chars_last,
      rematch009_in_chars        => Kernel_Nucleus_inst_rematch009_in_chars,
      rematch009_in_chars_count  => Kernel_Nucleus_inst_rematch009_in_chars_count,
      rematch009_in_unl_valid    => Kernel_Nucleus_inst_rematch009_in_unl_valid,
      rematch009_in_unl_ready    => Kernel_Nucleus_inst_rematch009_in_unl_ready,
      rematch009_in_unl_tag      => Kernel_Nucleus_inst_rematch009_in_unl_tag,
      rematch009_in_cmd_valid    => Kernel_Nucleus_inst_rematch009_in_cmd_valid,
      rematch009_in_cmd_ready    => Kernel_Nucleus_inst_rematch009_in_cmd_ready,
      rematch009_in_cmd_firstIdx => Kernel_Nucleus_inst_rematch009_in_cmd_firstIdx,
      rematch009_in_cmd_lastIdx  => Kernel_Nucleus_inst_rematch009_in_cmd_lastIdx,
      rematch009_in_cmd_ctrl     => Kernel_Nucleus_inst_rematch009_in_cmd_ctrl,
      rematch009_in_cmd_tag      => Kernel_Nucleus_inst_rematch009_in_cmd_tag,
      rematch010_in_valid        => Kernel_Nucleus_inst_rematch010_in_valid,
      rematch010_in_ready        => Kernel_Nucleus_inst_rematch010_in_ready,
      rematch010_in_dvalid       => Kernel_Nucleus_inst_rematch010_in_dvalid,
      rematch010_in_last         => Kernel_Nucleus_inst_rematch010_in_last,
      rematch010_in_length       => Kernel_Nucleus_inst_rematch010_in_length,
      rematch010_in_count        => Kernel_Nucleus_inst_rematch010_in_count,
      rematch010_in_chars_valid  => Kernel_Nucleus_inst_rematch010_in_chars_valid,
      rematch010_in_chars_ready  => Kernel_Nucleus_inst_rematch010_in_chars_ready,
      rematch010_in_chars_dvalid => Kernel_Nucleus_inst_rematch010_in_chars_dvalid,
      rematch010_in_chars_last   => Kernel_Nucleus_inst_rematch010_in_chars_last,
      rematch010_in_chars        => Kernel_Nucleus_inst_rematch010_in_chars,
      rematch010_in_chars_count  => Kernel_Nucleus_inst_rematch010_in_chars_count,
      rematch010_in_unl_valid    => Kernel_Nucleus_inst_rematch010_in_unl_valid,
      rematch010_in_unl_ready    => Kernel_Nucleus_inst_rematch010_in_unl_ready,
      rematch010_in_unl_tag      => Kernel_Nucleus_inst_rematch010_in_unl_tag,
      rematch010_in_cmd_valid    => Kernel_Nucleus_inst_rematch010_in_cmd_valid,
      rematch010_in_cmd_ready    => Kernel_Nucleus_inst_rematch010_in_cmd_ready,
      rematch010_in_cmd_firstIdx => Kernel_Nucleus_inst_rematch010_in_cmd_firstIdx,
      rematch010_in_cmd_lastIdx  => Kernel_Nucleus_inst_rematch010_in_cmd_lastIdx,
      rematch010_in_cmd_ctrl     => Kernel_Nucleus_inst_rematch010_in_cmd_ctrl,
      rematch010_in_cmd_tag      => Kernel_Nucleus_inst_rematch010_in_cmd_tag,
      rematch011_in_valid        => Kernel_Nucleus_inst_rematch011_in_valid,
      rematch011_in_ready        => Kernel_Nucleus_inst_rematch011_in_ready,
      rematch011_in_dvalid       => Kernel_Nucleus_inst_rematch011_in_dvalid,
      rematch011_in_last         => Kernel_Nucleus_inst_rematch011_in_last,
      rematch011_in_length       => Kernel_Nucleus_inst_rematch011_in_length,
      rematch011_in_count        => Kernel_Nucleus_inst_rematch011_in_count,
      rematch011_in_chars_valid  => Kernel_Nucleus_inst_rematch011_in_chars_valid,
      rematch011_in_chars_ready  => Kernel_Nucleus_inst_rematch011_in_chars_ready,
      rematch011_in_chars_dvalid => Kernel_Nucleus_inst_rematch011_in_chars_dvalid,
      rematch011_in_chars_last   => Kernel_Nucleus_inst_rematch011_in_chars_last,
      rematch011_in_chars        => Kernel_Nucleus_inst_rematch011_in_chars,
      rematch011_in_chars_count  => Kernel_Nucleus_inst_rematch011_in_chars_count,
      rematch011_in_unl_valid    => Kernel_Nucleus_inst_rematch011_in_unl_valid,
      rematch011_in_unl_ready    => Kernel_Nucleus_inst_rematch011_in_unl_ready,
      rematch011_in_unl_tag      => Kernel_Nucleus_inst_rematch011_in_unl_tag,
      rematch011_in_cmd_valid    => Kernel_Nucleus_inst_rematch011_in_cmd_valid,
      rematch011_in_cmd_ready    => Kernel_Nucleus_inst_rematch011_in_cmd_ready,
      rematch011_in_cmd_firstIdx => Kernel_Nucleus_inst_rematch011_in_cmd_firstIdx,
      rematch011_in_cmd_lastIdx  => Kernel_Nucleus_inst_rematch011_in_cmd_lastIdx,
      rematch011_in_cmd_ctrl     => Kernel_Nucleus_inst_rematch011_in_cmd_ctrl,
      rematch011_in_cmd_tag      => Kernel_Nucleus_inst_rematch011_in_cmd_tag,
      rematch012_in_valid        => Kernel_Nucleus_inst_rematch012_in_valid,
      rematch012_in_ready        => Kernel_Nucleus_inst_rematch012_in_ready,
      rematch012_in_dvalid       => Kernel_Nucleus_inst_rematch012_in_dvalid,
      rematch012_in_last         => Kernel_Nucleus_inst_rematch012_in_last,
      rematch012_in_length       => Kernel_Nucleus_inst_rematch012_in_length,
      rematch012_in_count        => Kernel_Nucleus_inst_rematch012_in_count,
      rematch012_in_chars_valid  => Kernel_Nucleus_inst_rematch012_in_chars_valid,
      rematch012_in_chars_ready  => Kernel_Nucleus_inst_rematch012_in_chars_ready,
      rematch012_in_chars_dvalid => Kernel_Nucleus_inst_rematch012_in_chars_dvalid,
      rematch012_in_chars_last   => Kernel_Nucleus_inst_rematch012_in_chars_last,
      rematch012_in_chars        => Kernel_Nucleus_inst_rematch012_in_chars,
      rematch012_in_chars_count  => Kernel_Nucleus_inst_rematch012_in_chars_count,
      rematch012_in_unl_valid    => Kernel_Nucleus_inst_rematch012_in_unl_valid,
      rematch012_in_unl_ready    => Kernel_Nucleus_inst_rematch012_in_unl_ready,
      rematch012_in_unl_tag      => Kernel_Nucleus_inst_rematch012_in_unl_tag,
      rematch012_in_cmd_valid    => Kernel_Nucleus_inst_rematch012_in_cmd_valid,
      rematch012_in_cmd_ready    => Kernel_Nucleus_inst_rematch012_in_cmd_ready,
      rematch012_in_cmd_firstIdx => Kernel_Nucleus_inst_rematch012_in_cmd_firstIdx,
      rematch012_in_cmd_lastIdx  => Kernel_Nucleus_inst_rematch012_in_cmd_lastIdx,
      rematch012_in_cmd_ctrl     => Kernel_Nucleus_inst_rematch012_in_cmd_ctrl,
      rematch012_in_cmd_tag      => Kernel_Nucleus_inst_rematch012_in_cmd_tag,
      rematch013_in_valid        => Kernel_Nucleus_inst_rematch013_in_valid,
      rematch013_in_ready        => Kernel_Nucleus_inst_rematch013_in_ready,
      rematch013_in_dvalid       => Kernel_Nucleus_inst_rematch013_in_dvalid,
      rematch013_in_last         => Kernel_Nucleus_inst_rematch013_in_last,
      rematch013_in_length       => Kernel_Nucleus_inst_rematch013_in_length,
      rematch013_in_count        => Kernel_Nucleus_inst_rematch013_in_count,
      rematch013_in_chars_valid  => Kernel_Nucleus_inst_rematch013_in_chars_valid,
      rematch013_in_chars_ready  => Kernel_Nucleus_inst_rematch013_in_chars_ready,
      rematch013_in_chars_dvalid => Kernel_Nucleus_inst_rematch013_in_chars_dvalid,
      rematch013_in_chars_last   => Kernel_Nucleus_inst_rematch013_in_chars_last,
      rematch013_in_chars        => Kernel_Nucleus_inst_rematch013_in_chars,
      rematch013_in_chars_count  => Kernel_Nucleus_inst_rematch013_in_chars_count,
      rematch013_in_unl_valid    => Kernel_Nucleus_inst_rematch013_in_unl_valid,
      rematch013_in_unl_ready    => Kernel_Nucleus_inst_rematch013_in_unl_ready,
      rematch013_in_unl_tag      => Kernel_Nucleus_inst_rematch013_in_unl_tag,
      rematch013_in_cmd_valid    => Kernel_Nucleus_inst_rematch013_in_cmd_valid,
      rematch013_in_cmd_ready    => Kernel_Nucleus_inst_rematch013_in_cmd_ready,
      rematch013_in_cmd_firstIdx => Kernel_Nucleus_inst_rematch013_in_cmd_firstIdx,
      rematch013_in_cmd_lastIdx  => Kernel_Nucleus_inst_rematch013_in_cmd_lastIdx,
      rematch013_in_cmd_ctrl     => Kernel_Nucleus_inst_rematch013_in_cmd_ctrl,
      rematch013_in_cmd_tag      => Kernel_Nucleus_inst_rematch013_in_cmd_tag,
      rematch014_in_valid        => Kernel_Nucleus_inst_rematch014_in_valid,
      rematch014_in_ready        => Kernel_Nucleus_inst_rematch014_in_ready,
      rematch014_in_dvalid       => Kernel_Nucleus_inst_rematch014_in_dvalid,
      rematch014_in_last         => Kernel_Nucleus_inst_rematch014_in_last,
      rematch014_in_length       => Kernel_Nucleus_inst_rematch014_in_length,
      rematch014_in_count        => Kernel_Nucleus_inst_rematch014_in_count,
      rematch014_in_chars_valid  => Kernel_Nucleus_inst_rematch014_in_chars_valid,
      rematch014_in_chars_ready  => Kernel_Nucleus_inst_rematch014_in_chars_ready,
      rematch014_in_chars_dvalid => Kernel_Nucleus_inst_rematch014_in_chars_dvalid,
      rematch014_in_chars_last   => Kernel_Nucleus_inst_rematch014_in_chars_last,
      rematch014_in_chars        => Kernel_Nucleus_inst_rematch014_in_chars,
      rematch014_in_chars_count  => Kernel_Nucleus_inst_rematch014_in_chars_count,
      rematch014_in_unl_valid    => Kernel_Nucleus_inst_rematch014_in_unl_valid,
      rematch014_in_unl_ready    => Kernel_Nucleus_inst_rematch014_in_unl_ready,
      rematch014_in_unl_tag      => Kernel_Nucleus_inst_rematch014_in_unl_tag,
      rematch014_in_cmd_valid    => Kernel_Nucleus_inst_rematch014_in_cmd_valid,
      rematch014_in_cmd_ready    => Kernel_Nucleus_inst_rematch014_in_cmd_ready,
      rematch014_in_cmd_firstIdx => Kernel_Nucleus_inst_rematch014_in_cmd_firstIdx,
      rematch014_in_cmd_lastIdx  => Kernel_Nucleus_inst_rematch014_in_cmd_lastIdx,
      rematch014_in_cmd_ctrl     => Kernel_Nucleus_inst_rematch014_in_cmd_ctrl,
      rematch014_in_cmd_tag      => Kernel_Nucleus_inst_rematch014_in_cmd_tag,
      rematch015_in_valid        => Kernel_Nucleus_inst_rematch015_in_valid,
      rematch015_in_ready        => Kernel_Nucleus_inst_rematch015_in_ready,
      rematch015_in_dvalid       => Kernel_Nucleus_inst_rematch015_in_dvalid,
      rematch015_in_last         => Kernel_Nucleus_inst_rematch015_in_last,
      rematch015_in_length       => Kernel_Nucleus_inst_rematch015_in_length,
      rematch015_in_count        => Kernel_Nucleus_inst_rematch015_in_count,
      rematch015_in_chars_valid  => Kernel_Nucleus_inst_rematch015_in_chars_valid,
      rematch015_in_chars_ready  => Kernel_Nucleus_inst_rematch015_in_chars_ready,
      rematch015_in_chars_dvalid => Kernel_Nucleus_inst_rematch015_in_chars_dvalid,
      rematch015_in_chars_last   => Kernel_Nucleus_inst_rematch015_in_chars_last,
      rematch015_in_chars        => Kernel_Nucleus_inst_rematch015_in_chars,
      rematch015_in_chars_count  => Kernel_Nucleus_inst_rematch015_in_chars_count,
      rematch015_in_unl_valid    => Kernel_Nucleus_inst_rematch015_in_unl_valid,
      rematch015_in_unl_ready    => Kernel_Nucleus_inst_rematch015_in_unl_ready,
      rematch015_in_unl_tag      => Kernel_Nucleus_inst_rematch015_in_unl_tag,
      rematch015_in_cmd_valid    => Kernel_Nucleus_inst_rematch015_in_cmd_valid,
      rematch015_in_cmd_ready    => Kernel_Nucleus_inst_rematch015_in_cmd_ready,
      rematch015_in_cmd_firstIdx => Kernel_Nucleus_inst_rematch015_in_cmd_firstIdx,
      rematch015_in_cmd_lastIdx  => Kernel_Nucleus_inst_rematch015_in_cmd_lastIdx,
      rematch015_in_cmd_ctrl     => Kernel_Nucleus_inst_rematch015_in_cmd_ctrl,
      rematch015_in_cmd_tag      => Kernel_Nucleus_inst_rematch015_in_cmd_tag
    );

  Kernel_rematch000_inst : Kernel_rematch000
    generic map (
      INDEX_WIDTH                      => INDEX_WIDTH,
      TAG_WIDTH                        => TAG_WIDTH,
      REMATCH000_IN_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
      REMATCH000_IN_BUS_DATA_WIDTH     => BUS_DATA_WIDTH,
      REMATCH000_IN_BUS_LEN_WIDTH      => BUS_LEN_WIDTH,
      REMATCH000_IN_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
      REMATCH000_IN_BUS_BURST_MAX_LEN  => BUS_BURST_MAX_LEN
    )
    port map (
      bcd_clk                      => bcd_clk,
      bcd_reset                    => bcd_reset,
      kcd_clk                      => kcd_clk,
      kcd_reset                    => kcd_reset,
      rematch000_in_valid          => Kernel_rematch000_inst_rematch000_in_valid,
      rematch000_in_ready          => Kernel_rematch000_inst_rematch000_in_ready,
      rematch000_in_dvalid         => Kernel_rematch000_inst_rematch000_in_dvalid,
      rematch000_in_last           => Kernel_rematch000_inst_rematch000_in_last,
      rematch000_in_length         => Kernel_rematch000_inst_rematch000_in_length,
      rematch000_in_count          => Kernel_rematch000_inst_rematch000_in_count,
      rematch000_in_chars_valid    => Kernel_rematch000_inst_rematch000_in_chars_valid,
      rematch000_in_chars_ready    => Kernel_rematch000_inst_rematch000_in_chars_ready,
      rematch000_in_chars_dvalid   => Kernel_rematch000_inst_rematch000_in_chars_dvalid,
      rematch000_in_chars_last     => Kernel_rematch000_inst_rematch000_in_chars_last,
      rematch000_in_chars          => Kernel_rematch000_inst_rematch000_in_chars,
      rematch000_in_chars_count    => Kernel_rematch000_inst_rematch000_in_chars_count,
      rematch000_in_bus_rreq_valid => Kernel_rematch000_inst_rematch000_in_bus_rreq_valid,
      rematch000_in_bus_rreq_ready => Kernel_rematch000_inst_rematch000_in_bus_rreq_ready,
      rematch000_in_bus_rreq_addr  => Kernel_rematch000_inst_rematch000_in_bus_rreq_addr,
      rematch000_in_bus_rreq_len   => Kernel_rematch000_inst_rematch000_in_bus_rreq_len,
      rematch000_in_bus_rdat_valid => Kernel_rematch000_inst_rematch000_in_bus_rdat_valid,
      rematch000_in_bus_rdat_ready => Kernel_rematch000_inst_rematch000_in_bus_rdat_ready,
      rematch000_in_bus_rdat_data  => Kernel_rematch000_inst_rematch000_in_bus_rdat_data,
      rematch000_in_bus_rdat_last  => Kernel_rematch000_inst_rematch000_in_bus_rdat_last,
      rematch000_in_cmd_valid      => Kernel_rematch000_inst_rematch000_in_cmd_valid,
      rematch000_in_cmd_ready      => Kernel_rematch000_inst_rematch000_in_cmd_ready,
      rematch000_in_cmd_firstIdx   => Kernel_rematch000_inst_rematch000_in_cmd_firstIdx,
      rematch000_in_cmd_lastIdx    => Kernel_rematch000_inst_rematch000_in_cmd_lastIdx,
      rematch000_in_cmd_ctrl       => Kernel_rematch000_inst_rematch000_in_cmd_ctrl,
      rematch000_in_cmd_tag        => Kernel_rematch000_inst_rematch000_in_cmd_tag,
      rematch000_in_unl_valid      => Kernel_rematch000_inst_rematch000_in_unl_valid,
      rematch000_in_unl_ready      => Kernel_rematch000_inst_rematch000_in_unl_ready,
      rematch000_in_unl_tag        => Kernel_rematch000_inst_rematch000_in_unl_tag
    );

  Kernel_rematch001_inst : Kernel_rematch001
    generic map (
      INDEX_WIDTH                      => INDEX_WIDTH,
      TAG_WIDTH                        => TAG_WIDTH,
      REMATCH001_IN_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
      REMATCH001_IN_BUS_DATA_WIDTH     => BUS_DATA_WIDTH,
      REMATCH001_IN_BUS_LEN_WIDTH      => BUS_LEN_WIDTH,
      REMATCH001_IN_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
      REMATCH001_IN_BUS_BURST_MAX_LEN  => BUS_BURST_MAX_LEN
    )
    port map (
      bcd_clk                      => bcd_clk,
      bcd_reset                    => bcd_reset,
      kcd_clk                      => kcd_clk,
      kcd_reset                    => kcd_reset,
      rematch001_in_valid          => Kernel_rematch001_inst_rematch001_in_valid,
      rematch001_in_ready          => Kernel_rematch001_inst_rematch001_in_ready,
      rematch001_in_dvalid         => Kernel_rematch001_inst_rematch001_in_dvalid,
      rematch001_in_last           => Kernel_rematch001_inst_rematch001_in_last,
      rematch001_in_length         => Kernel_rematch001_inst_rematch001_in_length,
      rematch001_in_count          => Kernel_rematch001_inst_rematch001_in_count,
      rematch001_in_chars_valid    => Kernel_rematch001_inst_rematch001_in_chars_valid,
      rematch001_in_chars_ready    => Kernel_rematch001_inst_rematch001_in_chars_ready,
      rematch001_in_chars_dvalid   => Kernel_rematch001_inst_rematch001_in_chars_dvalid,
      rematch001_in_chars_last     => Kernel_rematch001_inst_rematch001_in_chars_last,
      rematch001_in_chars          => Kernel_rematch001_inst_rematch001_in_chars,
      rematch001_in_chars_count    => Kernel_rematch001_inst_rematch001_in_chars_count,
      rematch001_in_bus_rreq_valid => Kernel_rematch001_inst_rematch001_in_bus_rreq_valid,
      rematch001_in_bus_rreq_ready => Kernel_rematch001_inst_rematch001_in_bus_rreq_ready,
      rematch001_in_bus_rreq_addr  => Kernel_rematch001_inst_rematch001_in_bus_rreq_addr,
      rematch001_in_bus_rreq_len   => Kernel_rematch001_inst_rematch001_in_bus_rreq_len,
      rematch001_in_bus_rdat_valid => Kernel_rematch001_inst_rematch001_in_bus_rdat_valid,
      rematch001_in_bus_rdat_ready => Kernel_rematch001_inst_rematch001_in_bus_rdat_ready,
      rematch001_in_bus_rdat_data  => Kernel_rematch001_inst_rematch001_in_bus_rdat_data,
      rematch001_in_bus_rdat_last  => Kernel_rematch001_inst_rematch001_in_bus_rdat_last,
      rematch001_in_cmd_valid      => Kernel_rematch001_inst_rematch001_in_cmd_valid,
      rematch001_in_cmd_ready      => Kernel_rematch001_inst_rematch001_in_cmd_ready,
      rematch001_in_cmd_firstIdx   => Kernel_rematch001_inst_rematch001_in_cmd_firstIdx,
      rematch001_in_cmd_lastIdx    => Kernel_rematch001_inst_rematch001_in_cmd_lastIdx,
      rematch001_in_cmd_ctrl       => Kernel_rematch001_inst_rematch001_in_cmd_ctrl,
      rematch001_in_cmd_tag        => Kernel_rematch001_inst_rematch001_in_cmd_tag,
      rematch001_in_unl_valid      => Kernel_rematch001_inst_rematch001_in_unl_valid,
      rematch001_in_unl_ready      => Kernel_rematch001_inst_rematch001_in_unl_ready,
      rematch001_in_unl_tag        => Kernel_rematch001_inst_rematch001_in_unl_tag
    );

  Kernel_rematch002_inst : Kernel_rematch002
    generic map (
      INDEX_WIDTH                      => INDEX_WIDTH,
      TAG_WIDTH                        => TAG_WIDTH,
      REMATCH002_IN_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
      REMATCH002_IN_BUS_DATA_WIDTH     => BUS_DATA_WIDTH,
      REMATCH002_IN_BUS_LEN_WIDTH      => BUS_LEN_WIDTH,
      REMATCH002_IN_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
      REMATCH002_IN_BUS_BURST_MAX_LEN  => BUS_BURST_MAX_LEN
    )
    port map (
      bcd_clk                      => bcd_clk,
      bcd_reset                    => bcd_reset,
      kcd_clk                      => kcd_clk,
      kcd_reset                    => kcd_reset,
      rematch002_in_valid          => Kernel_rematch002_inst_rematch002_in_valid,
      rematch002_in_ready          => Kernel_rematch002_inst_rematch002_in_ready,
      rematch002_in_dvalid         => Kernel_rematch002_inst_rematch002_in_dvalid,
      rematch002_in_last           => Kernel_rematch002_inst_rematch002_in_last,
      rematch002_in_length         => Kernel_rematch002_inst_rematch002_in_length,
      rematch002_in_count          => Kernel_rematch002_inst_rematch002_in_count,
      rematch002_in_chars_valid    => Kernel_rematch002_inst_rematch002_in_chars_valid,
      rematch002_in_chars_ready    => Kernel_rematch002_inst_rematch002_in_chars_ready,
      rematch002_in_chars_dvalid   => Kernel_rematch002_inst_rematch002_in_chars_dvalid,
      rematch002_in_chars_last     => Kernel_rematch002_inst_rematch002_in_chars_last,
      rematch002_in_chars          => Kernel_rematch002_inst_rematch002_in_chars,
      rematch002_in_chars_count    => Kernel_rematch002_inst_rematch002_in_chars_count,
      rematch002_in_bus_rreq_valid => Kernel_rematch002_inst_rematch002_in_bus_rreq_valid,
      rematch002_in_bus_rreq_ready => Kernel_rematch002_inst_rematch002_in_bus_rreq_ready,
      rematch002_in_bus_rreq_addr  => Kernel_rematch002_inst_rematch002_in_bus_rreq_addr,
      rematch002_in_bus_rreq_len   => Kernel_rematch002_inst_rematch002_in_bus_rreq_len,
      rematch002_in_bus_rdat_valid => Kernel_rematch002_inst_rematch002_in_bus_rdat_valid,
      rematch002_in_bus_rdat_ready => Kernel_rematch002_inst_rematch002_in_bus_rdat_ready,
      rematch002_in_bus_rdat_data  => Kernel_rematch002_inst_rematch002_in_bus_rdat_data,
      rematch002_in_bus_rdat_last  => Kernel_rematch002_inst_rematch002_in_bus_rdat_last,
      rematch002_in_cmd_valid      => Kernel_rematch002_inst_rematch002_in_cmd_valid,
      rematch002_in_cmd_ready      => Kernel_rematch002_inst_rematch002_in_cmd_ready,
      rematch002_in_cmd_firstIdx   => Kernel_rematch002_inst_rematch002_in_cmd_firstIdx,
      rematch002_in_cmd_lastIdx    => Kernel_rematch002_inst_rematch002_in_cmd_lastIdx,
      rematch002_in_cmd_ctrl       => Kernel_rematch002_inst_rematch002_in_cmd_ctrl,
      rematch002_in_cmd_tag        => Kernel_rematch002_inst_rematch002_in_cmd_tag,
      rematch002_in_unl_valid      => Kernel_rematch002_inst_rematch002_in_unl_valid,
      rematch002_in_unl_ready      => Kernel_rematch002_inst_rematch002_in_unl_ready,
      rematch002_in_unl_tag        => Kernel_rematch002_inst_rematch002_in_unl_tag
    );

  Kernel_rematch003_inst : Kernel_rematch003
    generic map (
      INDEX_WIDTH                      => INDEX_WIDTH,
      TAG_WIDTH                        => TAG_WIDTH,
      REMATCH003_IN_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
      REMATCH003_IN_BUS_DATA_WIDTH     => BUS_DATA_WIDTH,
      REMATCH003_IN_BUS_LEN_WIDTH      => BUS_LEN_WIDTH,
      REMATCH003_IN_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
      REMATCH003_IN_BUS_BURST_MAX_LEN  => BUS_BURST_MAX_LEN
    )
    port map (
      bcd_clk                      => bcd_clk,
      bcd_reset                    => bcd_reset,
      kcd_clk                      => kcd_clk,
      kcd_reset                    => kcd_reset,
      rematch003_in_valid          => Kernel_rematch003_inst_rematch003_in_valid,
      rematch003_in_ready          => Kernel_rematch003_inst_rematch003_in_ready,
      rematch003_in_dvalid         => Kernel_rematch003_inst_rematch003_in_dvalid,
      rematch003_in_last           => Kernel_rematch003_inst_rematch003_in_last,
      rematch003_in_length         => Kernel_rematch003_inst_rematch003_in_length,
      rematch003_in_count          => Kernel_rematch003_inst_rematch003_in_count,
      rematch003_in_chars_valid    => Kernel_rematch003_inst_rematch003_in_chars_valid,
      rematch003_in_chars_ready    => Kernel_rematch003_inst_rematch003_in_chars_ready,
      rematch003_in_chars_dvalid   => Kernel_rematch003_inst_rematch003_in_chars_dvalid,
      rematch003_in_chars_last     => Kernel_rematch003_inst_rematch003_in_chars_last,
      rematch003_in_chars          => Kernel_rematch003_inst_rematch003_in_chars,
      rematch003_in_chars_count    => Kernel_rematch003_inst_rematch003_in_chars_count,
      rematch003_in_bus_rreq_valid => Kernel_rematch003_inst_rematch003_in_bus_rreq_valid,
      rematch003_in_bus_rreq_ready => Kernel_rematch003_inst_rematch003_in_bus_rreq_ready,
      rematch003_in_bus_rreq_addr  => Kernel_rematch003_inst_rematch003_in_bus_rreq_addr,
      rematch003_in_bus_rreq_len   => Kernel_rematch003_inst_rematch003_in_bus_rreq_len,
      rematch003_in_bus_rdat_valid => Kernel_rematch003_inst_rematch003_in_bus_rdat_valid,
      rematch003_in_bus_rdat_ready => Kernel_rematch003_inst_rematch003_in_bus_rdat_ready,
      rematch003_in_bus_rdat_data  => Kernel_rematch003_inst_rematch003_in_bus_rdat_data,
      rematch003_in_bus_rdat_last  => Kernel_rematch003_inst_rematch003_in_bus_rdat_last,
      rematch003_in_cmd_valid      => Kernel_rematch003_inst_rematch003_in_cmd_valid,
      rematch003_in_cmd_ready      => Kernel_rematch003_inst_rematch003_in_cmd_ready,
      rematch003_in_cmd_firstIdx   => Kernel_rematch003_inst_rematch003_in_cmd_firstIdx,
      rematch003_in_cmd_lastIdx    => Kernel_rematch003_inst_rematch003_in_cmd_lastIdx,
      rematch003_in_cmd_ctrl       => Kernel_rematch003_inst_rematch003_in_cmd_ctrl,
      rematch003_in_cmd_tag        => Kernel_rematch003_inst_rematch003_in_cmd_tag,
      rematch003_in_unl_valid      => Kernel_rematch003_inst_rematch003_in_unl_valid,
      rematch003_in_unl_ready      => Kernel_rematch003_inst_rematch003_in_unl_ready,
      rematch003_in_unl_tag        => Kernel_rematch003_inst_rematch003_in_unl_tag
    );

  Kernel_rematch004_inst : Kernel_rematch004
    generic map (
      INDEX_WIDTH                      => INDEX_WIDTH,
      TAG_WIDTH                        => TAG_WIDTH,
      REMATCH004_IN_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
      REMATCH004_IN_BUS_DATA_WIDTH     => BUS_DATA_WIDTH,
      REMATCH004_IN_BUS_LEN_WIDTH      => BUS_LEN_WIDTH,
      REMATCH004_IN_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
      REMATCH004_IN_BUS_BURST_MAX_LEN  => BUS_BURST_MAX_LEN
    )
    port map (
      bcd_clk                      => bcd_clk,
      bcd_reset                    => bcd_reset,
      kcd_clk                      => kcd_clk,
      kcd_reset                    => kcd_reset,
      rematch004_in_valid          => Kernel_rematch004_inst_rematch004_in_valid,
      rematch004_in_ready          => Kernel_rematch004_inst_rematch004_in_ready,
      rematch004_in_dvalid         => Kernel_rematch004_inst_rematch004_in_dvalid,
      rematch004_in_last           => Kernel_rematch004_inst_rematch004_in_last,
      rematch004_in_length         => Kernel_rematch004_inst_rematch004_in_length,
      rematch004_in_count          => Kernel_rematch004_inst_rematch004_in_count,
      rematch004_in_chars_valid    => Kernel_rematch004_inst_rematch004_in_chars_valid,
      rematch004_in_chars_ready    => Kernel_rematch004_inst_rematch004_in_chars_ready,
      rematch004_in_chars_dvalid   => Kernel_rematch004_inst_rematch004_in_chars_dvalid,
      rematch004_in_chars_last     => Kernel_rematch004_inst_rematch004_in_chars_last,
      rematch004_in_chars          => Kernel_rematch004_inst_rematch004_in_chars,
      rematch004_in_chars_count    => Kernel_rematch004_inst_rematch004_in_chars_count,
      rematch004_in_bus_rreq_valid => Kernel_rematch004_inst_rematch004_in_bus_rreq_valid,
      rematch004_in_bus_rreq_ready => Kernel_rematch004_inst_rematch004_in_bus_rreq_ready,
      rematch004_in_bus_rreq_addr  => Kernel_rematch004_inst_rematch004_in_bus_rreq_addr,
      rematch004_in_bus_rreq_len   => Kernel_rematch004_inst_rematch004_in_bus_rreq_len,
      rematch004_in_bus_rdat_valid => Kernel_rematch004_inst_rematch004_in_bus_rdat_valid,
      rematch004_in_bus_rdat_ready => Kernel_rematch004_inst_rematch004_in_bus_rdat_ready,
      rematch004_in_bus_rdat_data  => Kernel_rematch004_inst_rematch004_in_bus_rdat_data,
      rematch004_in_bus_rdat_last  => Kernel_rematch004_inst_rematch004_in_bus_rdat_last,
      rematch004_in_cmd_valid      => Kernel_rematch004_inst_rematch004_in_cmd_valid,
      rematch004_in_cmd_ready      => Kernel_rematch004_inst_rematch004_in_cmd_ready,
      rematch004_in_cmd_firstIdx   => Kernel_rematch004_inst_rematch004_in_cmd_firstIdx,
      rematch004_in_cmd_lastIdx    => Kernel_rematch004_inst_rematch004_in_cmd_lastIdx,
      rematch004_in_cmd_ctrl       => Kernel_rematch004_inst_rematch004_in_cmd_ctrl,
      rematch004_in_cmd_tag        => Kernel_rematch004_inst_rematch004_in_cmd_tag,
      rematch004_in_unl_valid      => Kernel_rematch004_inst_rematch004_in_unl_valid,
      rematch004_in_unl_ready      => Kernel_rematch004_inst_rematch004_in_unl_ready,
      rematch004_in_unl_tag        => Kernel_rematch004_inst_rematch004_in_unl_tag
    );

  Kernel_rematch005_inst : Kernel_rematch005
    generic map (
      INDEX_WIDTH                      => INDEX_WIDTH,
      TAG_WIDTH                        => TAG_WIDTH,
      REMATCH005_IN_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
      REMATCH005_IN_BUS_DATA_WIDTH     => BUS_DATA_WIDTH,
      REMATCH005_IN_BUS_LEN_WIDTH      => BUS_LEN_WIDTH,
      REMATCH005_IN_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
      REMATCH005_IN_BUS_BURST_MAX_LEN  => BUS_BURST_MAX_LEN
    )
    port map (
      bcd_clk                      => bcd_clk,
      bcd_reset                    => bcd_reset,
      kcd_clk                      => kcd_clk,
      kcd_reset                    => kcd_reset,
      rematch005_in_valid          => Kernel_rematch005_inst_rematch005_in_valid,
      rematch005_in_ready          => Kernel_rematch005_inst_rematch005_in_ready,
      rematch005_in_dvalid         => Kernel_rematch005_inst_rematch005_in_dvalid,
      rematch005_in_last           => Kernel_rematch005_inst_rematch005_in_last,
      rematch005_in_length         => Kernel_rematch005_inst_rematch005_in_length,
      rematch005_in_count          => Kernel_rematch005_inst_rematch005_in_count,
      rematch005_in_chars_valid    => Kernel_rematch005_inst_rematch005_in_chars_valid,
      rematch005_in_chars_ready    => Kernel_rematch005_inst_rematch005_in_chars_ready,
      rematch005_in_chars_dvalid   => Kernel_rematch005_inst_rematch005_in_chars_dvalid,
      rematch005_in_chars_last     => Kernel_rematch005_inst_rematch005_in_chars_last,
      rematch005_in_chars          => Kernel_rematch005_inst_rematch005_in_chars,
      rematch005_in_chars_count    => Kernel_rematch005_inst_rematch005_in_chars_count,
      rematch005_in_bus_rreq_valid => Kernel_rematch005_inst_rematch005_in_bus_rreq_valid,
      rematch005_in_bus_rreq_ready => Kernel_rematch005_inst_rematch005_in_bus_rreq_ready,
      rematch005_in_bus_rreq_addr  => Kernel_rematch005_inst_rematch005_in_bus_rreq_addr,
      rematch005_in_bus_rreq_len   => Kernel_rematch005_inst_rematch005_in_bus_rreq_len,
      rematch005_in_bus_rdat_valid => Kernel_rematch005_inst_rematch005_in_bus_rdat_valid,
      rematch005_in_bus_rdat_ready => Kernel_rematch005_inst_rematch005_in_bus_rdat_ready,
      rematch005_in_bus_rdat_data  => Kernel_rematch005_inst_rematch005_in_bus_rdat_data,
      rematch005_in_bus_rdat_last  => Kernel_rematch005_inst_rematch005_in_bus_rdat_last,
      rematch005_in_cmd_valid      => Kernel_rematch005_inst_rematch005_in_cmd_valid,
      rematch005_in_cmd_ready      => Kernel_rematch005_inst_rematch005_in_cmd_ready,
      rematch005_in_cmd_firstIdx   => Kernel_rematch005_inst_rematch005_in_cmd_firstIdx,
      rematch005_in_cmd_lastIdx    => Kernel_rematch005_inst_rematch005_in_cmd_lastIdx,
      rematch005_in_cmd_ctrl       => Kernel_rematch005_inst_rematch005_in_cmd_ctrl,
      rematch005_in_cmd_tag        => Kernel_rematch005_inst_rematch005_in_cmd_tag,
      rematch005_in_unl_valid      => Kernel_rematch005_inst_rematch005_in_unl_valid,
      rematch005_in_unl_ready      => Kernel_rematch005_inst_rematch005_in_unl_ready,
      rematch005_in_unl_tag        => Kernel_rematch005_inst_rematch005_in_unl_tag
    );

  Kernel_rematch006_inst : Kernel_rematch006
    generic map (
      INDEX_WIDTH                      => INDEX_WIDTH,
      TAG_WIDTH                        => TAG_WIDTH,
      REMATCH006_IN_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
      REMATCH006_IN_BUS_DATA_WIDTH     => BUS_DATA_WIDTH,
      REMATCH006_IN_BUS_LEN_WIDTH      => BUS_LEN_WIDTH,
      REMATCH006_IN_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
      REMATCH006_IN_BUS_BURST_MAX_LEN  => BUS_BURST_MAX_LEN
    )
    port map (
      bcd_clk                      => bcd_clk,
      bcd_reset                    => bcd_reset,
      kcd_clk                      => kcd_clk,
      kcd_reset                    => kcd_reset,
      rematch006_in_valid          => Kernel_rematch006_inst_rematch006_in_valid,
      rematch006_in_ready          => Kernel_rematch006_inst_rematch006_in_ready,
      rematch006_in_dvalid         => Kernel_rematch006_inst_rematch006_in_dvalid,
      rematch006_in_last           => Kernel_rematch006_inst_rematch006_in_last,
      rematch006_in_length         => Kernel_rematch006_inst_rematch006_in_length,
      rematch006_in_count          => Kernel_rematch006_inst_rematch006_in_count,
      rematch006_in_chars_valid    => Kernel_rematch006_inst_rematch006_in_chars_valid,
      rematch006_in_chars_ready    => Kernel_rematch006_inst_rematch006_in_chars_ready,
      rematch006_in_chars_dvalid   => Kernel_rematch006_inst_rematch006_in_chars_dvalid,
      rematch006_in_chars_last     => Kernel_rematch006_inst_rematch006_in_chars_last,
      rematch006_in_chars          => Kernel_rematch006_inst_rematch006_in_chars,
      rematch006_in_chars_count    => Kernel_rematch006_inst_rematch006_in_chars_count,
      rematch006_in_bus_rreq_valid => Kernel_rematch006_inst_rematch006_in_bus_rreq_valid,
      rematch006_in_bus_rreq_ready => Kernel_rematch006_inst_rematch006_in_bus_rreq_ready,
      rematch006_in_bus_rreq_addr  => Kernel_rematch006_inst_rematch006_in_bus_rreq_addr,
      rematch006_in_bus_rreq_len   => Kernel_rematch006_inst_rematch006_in_bus_rreq_len,
      rematch006_in_bus_rdat_valid => Kernel_rematch006_inst_rematch006_in_bus_rdat_valid,
      rematch006_in_bus_rdat_ready => Kernel_rematch006_inst_rematch006_in_bus_rdat_ready,
      rematch006_in_bus_rdat_data  => Kernel_rematch006_inst_rematch006_in_bus_rdat_data,
      rematch006_in_bus_rdat_last  => Kernel_rematch006_inst_rematch006_in_bus_rdat_last,
      rematch006_in_cmd_valid      => Kernel_rematch006_inst_rematch006_in_cmd_valid,
      rematch006_in_cmd_ready      => Kernel_rematch006_inst_rematch006_in_cmd_ready,
      rematch006_in_cmd_firstIdx   => Kernel_rematch006_inst_rematch006_in_cmd_firstIdx,
      rematch006_in_cmd_lastIdx    => Kernel_rematch006_inst_rematch006_in_cmd_lastIdx,
      rematch006_in_cmd_ctrl       => Kernel_rematch006_inst_rematch006_in_cmd_ctrl,
      rematch006_in_cmd_tag        => Kernel_rematch006_inst_rematch006_in_cmd_tag,
      rematch006_in_unl_valid      => Kernel_rematch006_inst_rematch006_in_unl_valid,
      rematch006_in_unl_ready      => Kernel_rematch006_inst_rematch006_in_unl_ready,
      rematch006_in_unl_tag        => Kernel_rematch006_inst_rematch006_in_unl_tag
    );

  Kernel_rematch007_inst : Kernel_rematch007
    generic map (
      INDEX_WIDTH                      => INDEX_WIDTH,
      TAG_WIDTH                        => TAG_WIDTH,
      REMATCH007_IN_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
      REMATCH007_IN_BUS_DATA_WIDTH     => BUS_DATA_WIDTH,
      REMATCH007_IN_BUS_LEN_WIDTH      => BUS_LEN_WIDTH,
      REMATCH007_IN_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
      REMATCH007_IN_BUS_BURST_MAX_LEN  => BUS_BURST_MAX_LEN
    )
    port map (
      bcd_clk                      => bcd_clk,
      bcd_reset                    => bcd_reset,
      kcd_clk                      => kcd_clk,
      kcd_reset                    => kcd_reset,
      rematch007_in_valid          => Kernel_rematch007_inst_rematch007_in_valid,
      rematch007_in_ready          => Kernel_rematch007_inst_rematch007_in_ready,
      rematch007_in_dvalid         => Kernel_rematch007_inst_rematch007_in_dvalid,
      rematch007_in_last           => Kernel_rematch007_inst_rematch007_in_last,
      rematch007_in_length         => Kernel_rematch007_inst_rematch007_in_length,
      rematch007_in_count          => Kernel_rematch007_inst_rematch007_in_count,
      rematch007_in_chars_valid    => Kernel_rematch007_inst_rematch007_in_chars_valid,
      rematch007_in_chars_ready    => Kernel_rematch007_inst_rematch007_in_chars_ready,
      rematch007_in_chars_dvalid   => Kernel_rematch007_inst_rematch007_in_chars_dvalid,
      rematch007_in_chars_last     => Kernel_rematch007_inst_rematch007_in_chars_last,
      rematch007_in_chars          => Kernel_rematch007_inst_rematch007_in_chars,
      rematch007_in_chars_count    => Kernel_rematch007_inst_rematch007_in_chars_count,
      rematch007_in_bus_rreq_valid => Kernel_rematch007_inst_rematch007_in_bus_rreq_valid,
      rematch007_in_bus_rreq_ready => Kernel_rematch007_inst_rematch007_in_bus_rreq_ready,
      rematch007_in_bus_rreq_addr  => Kernel_rematch007_inst_rematch007_in_bus_rreq_addr,
      rematch007_in_bus_rreq_len   => Kernel_rematch007_inst_rematch007_in_bus_rreq_len,
      rematch007_in_bus_rdat_valid => Kernel_rematch007_inst_rematch007_in_bus_rdat_valid,
      rematch007_in_bus_rdat_ready => Kernel_rematch007_inst_rematch007_in_bus_rdat_ready,
      rematch007_in_bus_rdat_data  => Kernel_rematch007_inst_rematch007_in_bus_rdat_data,
      rematch007_in_bus_rdat_last  => Kernel_rematch007_inst_rematch007_in_bus_rdat_last,
      rematch007_in_cmd_valid      => Kernel_rematch007_inst_rematch007_in_cmd_valid,
      rematch007_in_cmd_ready      => Kernel_rematch007_inst_rematch007_in_cmd_ready,
      rematch007_in_cmd_firstIdx   => Kernel_rematch007_inst_rematch007_in_cmd_firstIdx,
      rematch007_in_cmd_lastIdx    => Kernel_rematch007_inst_rematch007_in_cmd_lastIdx,
      rematch007_in_cmd_ctrl       => Kernel_rematch007_inst_rematch007_in_cmd_ctrl,
      rematch007_in_cmd_tag        => Kernel_rematch007_inst_rematch007_in_cmd_tag,
      rematch007_in_unl_valid      => Kernel_rematch007_inst_rematch007_in_unl_valid,
      rematch007_in_unl_ready      => Kernel_rematch007_inst_rematch007_in_unl_ready,
      rematch007_in_unl_tag        => Kernel_rematch007_inst_rematch007_in_unl_tag
    );

  Kernel_rematch008_inst : Kernel_rematch008
    generic map (
      INDEX_WIDTH                      => INDEX_WIDTH,
      TAG_WIDTH                        => TAG_WIDTH,
      REMATCH008_IN_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
      REMATCH008_IN_BUS_DATA_WIDTH     => BUS_DATA_WIDTH,
      REMATCH008_IN_BUS_LEN_WIDTH      => BUS_LEN_WIDTH,
      REMATCH008_IN_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
      REMATCH008_IN_BUS_BURST_MAX_LEN  => BUS_BURST_MAX_LEN
    )
    port map (
      bcd_clk                      => bcd_clk,
      bcd_reset                    => bcd_reset,
      kcd_clk                      => kcd_clk,
      kcd_reset                    => kcd_reset,
      rematch008_in_valid          => Kernel_rematch008_inst_rematch008_in_valid,
      rematch008_in_ready          => Kernel_rematch008_inst_rematch008_in_ready,
      rematch008_in_dvalid         => Kernel_rematch008_inst_rematch008_in_dvalid,
      rematch008_in_last           => Kernel_rematch008_inst_rematch008_in_last,
      rematch008_in_length         => Kernel_rematch008_inst_rematch008_in_length,
      rematch008_in_count          => Kernel_rematch008_inst_rematch008_in_count,
      rematch008_in_chars_valid    => Kernel_rematch008_inst_rematch008_in_chars_valid,
      rematch008_in_chars_ready    => Kernel_rematch008_inst_rematch008_in_chars_ready,
      rematch008_in_chars_dvalid   => Kernel_rematch008_inst_rematch008_in_chars_dvalid,
      rematch008_in_chars_last     => Kernel_rematch008_inst_rematch008_in_chars_last,
      rematch008_in_chars          => Kernel_rematch008_inst_rematch008_in_chars,
      rematch008_in_chars_count    => Kernel_rematch008_inst_rematch008_in_chars_count,
      rematch008_in_bus_rreq_valid => Kernel_rematch008_inst_rematch008_in_bus_rreq_valid,
      rematch008_in_bus_rreq_ready => Kernel_rematch008_inst_rematch008_in_bus_rreq_ready,
      rematch008_in_bus_rreq_addr  => Kernel_rematch008_inst_rematch008_in_bus_rreq_addr,
      rematch008_in_bus_rreq_len   => Kernel_rematch008_inst_rematch008_in_bus_rreq_len,
      rematch008_in_bus_rdat_valid => Kernel_rematch008_inst_rematch008_in_bus_rdat_valid,
      rematch008_in_bus_rdat_ready => Kernel_rematch008_inst_rematch008_in_bus_rdat_ready,
      rematch008_in_bus_rdat_data  => Kernel_rematch008_inst_rematch008_in_bus_rdat_data,
      rematch008_in_bus_rdat_last  => Kernel_rematch008_inst_rematch008_in_bus_rdat_last,
      rematch008_in_cmd_valid      => Kernel_rematch008_inst_rematch008_in_cmd_valid,
      rematch008_in_cmd_ready      => Kernel_rematch008_inst_rematch008_in_cmd_ready,
      rematch008_in_cmd_firstIdx   => Kernel_rematch008_inst_rematch008_in_cmd_firstIdx,
      rematch008_in_cmd_lastIdx    => Kernel_rematch008_inst_rematch008_in_cmd_lastIdx,
      rematch008_in_cmd_ctrl       => Kernel_rematch008_inst_rematch008_in_cmd_ctrl,
      rematch008_in_cmd_tag        => Kernel_rematch008_inst_rematch008_in_cmd_tag,
      rematch008_in_unl_valid      => Kernel_rematch008_inst_rematch008_in_unl_valid,
      rematch008_in_unl_ready      => Kernel_rematch008_inst_rematch008_in_unl_ready,
      rematch008_in_unl_tag        => Kernel_rematch008_inst_rematch008_in_unl_tag
    );

  Kernel_rematch009_inst : Kernel_rematch009
    generic map (
      INDEX_WIDTH                      => INDEX_WIDTH,
      TAG_WIDTH                        => TAG_WIDTH,
      REMATCH009_IN_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
      REMATCH009_IN_BUS_DATA_WIDTH     => BUS_DATA_WIDTH,
      REMATCH009_IN_BUS_LEN_WIDTH      => BUS_LEN_WIDTH,
      REMATCH009_IN_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
      REMATCH009_IN_BUS_BURST_MAX_LEN  => BUS_BURST_MAX_LEN
    )
    port map (
      bcd_clk                      => bcd_clk,
      bcd_reset                    => bcd_reset,
      kcd_clk                      => kcd_clk,
      kcd_reset                    => kcd_reset,
      rematch009_in_valid          => Kernel_rematch009_inst_rematch009_in_valid,
      rematch009_in_ready          => Kernel_rematch009_inst_rematch009_in_ready,
      rematch009_in_dvalid         => Kernel_rematch009_inst_rematch009_in_dvalid,
      rematch009_in_last           => Kernel_rematch009_inst_rematch009_in_last,
      rematch009_in_length         => Kernel_rematch009_inst_rematch009_in_length,
      rematch009_in_count          => Kernel_rematch009_inst_rematch009_in_count,
      rematch009_in_chars_valid    => Kernel_rematch009_inst_rematch009_in_chars_valid,
      rematch009_in_chars_ready    => Kernel_rematch009_inst_rematch009_in_chars_ready,
      rematch009_in_chars_dvalid   => Kernel_rematch009_inst_rematch009_in_chars_dvalid,
      rematch009_in_chars_last     => Kernel_rematch009_inst_rematch009_in_chars_last,
      rematch009_in_chars          => Kernel_rematch009_inst_rematch009_in_chars,
      rematch009_in_chars_count    => Kernel_rematch009_inst_rematch009_in_chars_count,
      rematch009_in_bus_rreq_valid => Kernel_rematch009_inst_rematch009_in_bus_rreq_valid,
      rematch009_in_bus_rreq_ready => Kernel_rematch009_inst_rematch009_in_bus_rreq_ready,
      rematch009_in_bus_rreq_addr  => Kernel_rematch009_inst_rematch009_in_bus_rreq_addr,
      rematch009_in_bus_rreq_len   => Kernel_rematch009_inst_rematch009_in_bus_rreq_len,
      rematch009_in_bus_rdat_valid => Kernel_rematch009_inst_rematch009_in_bus_rdat_valid,
      rematch009_in_bus_rdat_ready => Kernel_rematch009_inst_rematch009_in_bus_rdat_ready,
      rematch009_in_bus_rdat_data  => Kernel_rematch009_inst_rematch009_in_bus_rdat_data,
      rematch009_in_bus_rdat_last  => Kernel_rematch009_inst_rematch009_in_bus_rdat_last,
      rematch009_in_cmd_valid      => Kernel_rematch009_inst_rematch009_in_cmd_valid,
      rematch009_in_cmd_ready      => Kernel_rematch009_inst_rematch009_in_cmd_ready,
      rematch009_in_cmd_firstIdx   => Kernel_rematch009_inst_rematch009_in_cmd_firstIdx,
      rematch009_in_cmd_lastIdx    => Kernel_rematch009_inst_rematch009_in_cmd_lastIdx,
      rematch009_in_cmd_ctrl       => Kernel_rematch009_inst_rematch009_in_cmd_ctrl,
      rematch009_in_cmd_tag        => Kernel_rematch009_inst_rematch009_in_cmd_tag,
      rematch009_in_unl_valid      => Kernel_rematch009_inst_rematch009_in_unl_valid,
      rematch009_in_unl_ready      => Kernel_rematch009_inst_rematch009_in_unl_ready,
      rematch009_in_unl_tag        => Kernel_rematch009_inst_rematch009_in_unl_tag
    );

  Kernel_rematch010_inst : Kernel_rematch010
    generic map (
      INDEX_WIDTH                      => INDEX_WIDTH,
      TAG_WIDTH                        => TAG_WIDTH,
      REMATCH010_IN_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
      REMATCH010_IN_BUS_DATA_WIDTH     => BUS_DATA_WIDTH,
      REMATCH010_IN_BUS_LEN_WIDTH      => BUS_LEN_WIDTH,
      REMATCH010_IN_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
      REMATCH010_IN_BUS_BURST_MAX_LEN  => BUS_BURST_MAX_LEN
    )
    port map (
      bcd_clk                      => bcd_clk,
      bcd_reset                    => bcd_reset,
      kcd_clk                      => kcd_clk,
      kcd_reset                    => kcd_reset,
      rematch010_in_valid          => Kernel_rematch010_inst_rematch010_in_valid,
      rematch010_in_ready          => Kernel_rematch010_inst_rematch010_in_ready,
      rematch010_in_dvalid         => Kernel_rematch010_inst_rematch010_in_dvalid,
      rematch010_in_last           => Kernel_rematch010_inst_rematch010_in_last,
      rematch010_in_length         => Kernel_rematch010_inst_rematch010_in_length,
      rematch010_in_count          => Kernel_rematch010_inst_rematch010_in_count,
      rematch010_in_chars_valid    => Kernel_rematch010_inst_rematch010_in_chars_valid,
      rematch010_in_chars_ready    => Kernel_rematch010_inst_rematch010_in_chars_ready,
      rematch010_in_chars_dvalid   => Kernel_rematch010_inst_rematch010_in_chars_dvalid,
      rematch010_in_chars_last     => Kernel_rematch010_inst_rematch010_in_chars_last,
      rematch010_in_chars          => Kernel_rematch010_inst_rematch010_in_chars,
      rematch010_in_chars_count    => Kernel_rematch010_inst_rematch010_in_chars_count,
      rematch010_in_bus_rreq_valid => Kernel_rematch010_inst_rematch010_in_bus_rreq_valid,
      rematch010_in_bus_rreq_ready => Kernel_rematch010_inst_rematch010_in_bus_rreq_ready,
      rematch010_in_bus_rreq_addr  => Kernel_rematch010_inst_rematch010_in_bus_rreq_addr,
      rematch010_in_bus_rreq_len   => Kernel_rematch010_inst_rematch010_in_bus_rreq_len,
      rematch010_in_bus_rdat_valid => Kernel_rematch010_inst_rematch010_in_bus_rdat_valid,
      rematch010_in_bus_rdat_ready => Kernel_rematch010_inst_rematch010_in_bus_rdat_ready,
      rematch010_in_bus_rdat_data  => Kernel_rematch010_inst_rematch010_in_bus_rdat_data,
      rematch010_in_bus_rdat_last  => Kernel_rematch010_inst_rematch010_in_bus_rdat_last,
      rematch010_in_cmd_valid      => Kernel_rematch010_inst_rematch010_in_cmd_valid,
      rematch010_in_cmd_ready      => Kernel_rematch010_inst_rematch010_in_cmd_ready,
      rematch010_in_cmd_firstIdx   => Kernel_rematch010_inst_rematch010_in_cmd_firstIdx,
      rematch010_in_cmd_lastIdx    => Kernel_rematch010_inst_rematch010_in_cmd_lastIdx,
      rematch010_in_cmd_ctrl       => Kernel_rematch010_inst_rematch010_in_cmd_ctrl,
      rematch010_in_cmd_tag        => Kernel_rematch010_inst_rematch010_in_cmd_tag,
      rematch010_in_unl_valid      => Kernel_rematch010_inst_rematch010_in_unl_valid,
      rematch010_in_unl_ready      => Kernel_rematch010_inst_rematch010_in_unl_ready,
      rematch010_in_unl_tag        => Kernel_rematch010_inst_rematch010_in_unl_tag
    );

  Kernel_rematch011_inst : Kernel_rematch011
    generic map (
      INDEX_WIDTH                      => INDEX_WIDTH,
      TAG_WIDTH                        => TAG_WIDTH,
      REMATCH011_IN_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
      REMATCH011_IN_BUS_DATA_WIDTH     => BUS_DATA_WIDTH,
      REMATCH011_IN_BUS_LEN_WIDTH      => BUS_LEN_WIDTH,
      REMATCH011_IN_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
      REMATCH011_IN_BUS_BURST_MAX_LEN  => BUS_BURST_MAX_LEN
    )
    port map (
      bcd_clk                      => bcd_clk,
      bcd_reset                    => bcd_reset,
      kcd_clk                      => kcd_clk,
      kcd_reset                    => kcd_reset,
      rematch011_in_valid          => Kernel_rematch011_inst_rematch011_in_valid,
      rematch011_in_ready          => Kernel_rematch011_inst_rematch011_in_ready,
      rematch011_in_dvalid         => Kernel_rematch011_inst_rematch011_in_dvalid,
      rematch011_in_last           => Kernel_rematch011_inst_rematch011_in_last,
      rematch011_in_length         => Kernel_rematch011_inst_rematch011_in_length,
      rematch011_in_count          => Kernel_rematch011_inst_rematch011_in_count,
      rematch011_in_chars_valid    => Kernel_rematch011_inst_rematch011_in_chars_valid,
      rematch011_in_chars_ready    => Kernel_rematch011_inst_rematch011_in_chars_ready,
      rematch011_in_chars_dvalid   => Kernel_rematch011_inst_rematch011_in_chars_dvalid,
      rematch011_in_chars_last     => Kernel_rematch011_inst_rematch011_in_chars_last,
      rematch011_in_chars          => Kernel_rematch011_inst_rematch011_in_chars,
      rematch011_in_chars_count    => Kernel_rematch011_inst_rematch011_in_chars_count,
      rematch011_in_bus_rreq_valid => Kernel_rematch011_inst_rematch011_in_bus_rreq_valid,
      rematch011_in_bus_rreq_ready => Kernel_rematch011_inst_rematch011_in_bus_rreq_ready,
      rematch011_in_bus_rreq_addr  => Kernel_rematch011_inst_rematch011_in_bus_rreq_addr,
      rematch011_in_bus_rreq_len   => Kernel_rematch011_inst_rematch011_in_bus_rreq_len,
      rematch011_in_bus_rdat_valid => Kernel_rematch011_inst_rematch011_in_bus_rdat_valid,
      rematch011_in_bus_rdat_ready => Kernel_rematch011_inst_rematch011_in_bus_rdat_ready,
      rematch011_in_bus_rdat_data  => Kernel_rematch011_inst_rematch011_in_bus_rdat_data,
      rematch011_in_bus_rdat_last  => Kernel_rematch011_inst_rematch011_in_bus_rdat_last,
      rematch011_in_cmd_valid      => Kernel_rematch011_inst_rematch011_in_cmd_valid,
      rematch011_in_cmd_ready      => Kernel_rematch011_inst_rematch011_in_cmd_ready,
      rematch011_in_cmd_firstIdx   => Kernel_rematch011_inst_rematch011_in_cmd_firstIdx,
      rematch011_in_cmd_lastIdx    => Kernel_rematch011_inst_rematch011_in_cmd_lastIdx,
      rematch011_in_cmd_ctrl       => Kernel_rematch011_inst_rematch011_in_cmd_ctrl,
      rematch011_in_cmd_tag        => Kernel_rematch011_inst_rematch011_in_cmd_tag,
      rematch011_in_unl_valid      => Kernel_rematch011_inst_rematch011_in_unl_valid,
      rematch011_in_unl_ready      => Kernel_rematch011_inst_rematch011_in_unl_ready,
      rematch011_in_unl_tag        => Kernel_rematch011_inst_rematch011_in_unl_tag
    );

  Kernel_rematch012_inst : Kernel_rematch012
    generic map (
      INDEX_WIDTH                      => INDEX_WIDTH,
      TAG_WIDTH                        => TAG_WIDTH,
      REMATCH012_IN_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
      REMATCH012_IN_BUS_DATA_WIDTH     => BUS_DATA_WIDTH,
      REMATCH012_IN_BUS_LEN_WIDTH      => BUS_LEN_WIDTH,
      REMATCH012_IN_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
      REMATCH012_IN_BUS_BURST_MAX_LEN  => BUS_BURST_MAX_LEN
    )
    port map (
      bcd_clk                      => bcd_clk,
      bcd_reset                    => bcd_reset,
      kcd_clk                      => kcd_clk,
      kcd_reset                    => kcd_reset,
      rematch012_in_valid          => Kernel_rematch012_inst_rematch012_in_valid,
      rematch012_in_ready          => Kernel_rematch012_inst_rematch012_in_ready,
      rematch012_in_dvalid         => Kernel_rematch012_inst_rematch012_in_dvalid,
      rematch012_in_last           => Kernel_rematch012_inst_rematch012_in_last,
      rematch012_in_length         => Kernel_rematch012_inst_rematch012_in_length,
      rematch012_in_count          => Kernel_rematch012_inst_rematch012_in_count,
      rematch012_in_chars_valid    => Kernel_rematch012_inst_rematch012_in_chars_valid,
      rematch012_in_chars_ready    => Kernel_rematch012_inst_rematch012_in_chars_ready,
      rematch012_in_chars_dvalid   => Kernel_rematch012_inst_rematch012_in_chars_dvalid,
      rematch012_in_chars_last     => Kernel_rematch012_inst_rematch012_in_chars_last,
      rematch012_in_chars          => Kernel_rematch012_inst_rematch012_in_chars,
      rematch012_in_chars_count    => Kernel_rematch012_inst_rematch012_in_chars_count,
      rematch012_in_bus_rreq_valid => Kernel_rematch012_inst_rematch012_in_bus_rreq_valid,
      rematch012_in_bus_rreq_ready => Kernel_rematch012_inst_rematch012_in_bus_rreq_ready,
      rematch012_in_bus_rreq_addr  => Kernel_rematch012_inst_rematch012_in_bus_rreq_addr,
      rematch012_in_bus_rreq_len   => Kernel_rematch012_inst_rematch012_in_bus_rreq_len,
      rematch012_in_bus_rdat_valid => Kernel_rematch012_inst_rematch012_in_bus_rdat_valid,
      rematch012_in_bus_rdat_ready => Kernel_rematch012_inst_rematch012_in_bus_rdat_ready,
      rematch012_in_bus_rdat_data  => Kernel_rematch012_inst_rematch012_in_bus_rdat_data,
      rematch012_in_bus_rdat_last  => Kernel_rematch012_inst_rematch012_in_bus_rdat_last,
      rematch012_in_cmd_valid      => Kernel_rematch012_inst_rematch012_in_cmd_valid,
      rematch012_in_cmd_ready      => Kernel_rematch012_inst_rematch012_in_cmd_ready,
      rematch012_in_cmd_firstIdx   => Kernel_rematch012_inst_rematch012_in_cmd_firstIdx,
      rematch012_in_cmd_lastIdx    => Kernel_rematch012_inst_rematch012_in_cmd_lastIdx,
      rematch012_in_cmd_ctrl       => Kernel_rematch012_inst_rematch012_in_cmd_ctrl,
      rematch012_in_cmd_tag        => Kernel_rematch012_inst_rematch012_in_cmd_tag,
      rematch012_in_unl_valid      => Kernel_rematch012_inst_rematch012_in_unl_valid,
      rematch012_in_unl_ready      => Kernel_rematch012_inst_rematch012_in_unl_ready,
      rematch012_in_unl_tag        => Kernel_rematch012_inst_rematch012_in_unl_tag
    );

  Kernel_rematch013_inst : Kernel_rematch013
    generic map (
      INDEX_WIDTH                      => INDEX_WIDTH,
      TAG_WIDTH                        => TAG_WIDTH,
      REMATCH013_IN_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
      REMATCH013_IN_BUS_DATA_WIDTH     => BUS_DATA_WIDTH,
      REMATCH013_IN_BUS_LEN_WIDTH      => BUS_LEN_WIDTH,
      REMATCH013_IN_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
      REMATCH013_IN_BUS_BURST_MAX_LEN  => BUS_BURST_MAX_LEN
    )
    port map (
      bcd_clk                      => bcd_clk,
      bcd_reset                    => bcd_reset,
      kcd_clk                      => kcd_clk,
      kcd_reset                    => kcd_reset,
      rematch013_in_valid          => Kernel_rematch013_inst_rematch013_in_valid,
      rematch013_in_ready          => Kernel_rematch013_inst_rematch013_in_ready,
      rematch013_in_dvalid         => Kernel_rematch013_inst_rematch013_in_dvalid,
      rematch013_in_last           => Kernel_rematch013_inst_rematch013_in_last,
      rematch013_in_length         => Kernel_rematch013_inst_rematch013_in_length,
      rematch013_in_count          => Kernel_rematch013_inst_rematch013_in_count,
      rematch013_in_chars_valid    => Kernel_rematch013_inst_rematch013_in_chars_valid,
      rematch013_in_chars_ready    => Kernel_rematch013_inst_rematch013_in_chars_ready,
      rematch013_in_chars_dvalid   => Kernel_rematch013_inst_rematch013_in_chars_dvalid,
      rematch013_in_chars_last     => Kernel_rematch013_inst_rematch013_in_chars_last,
      rematch013_in_chars          => Kernel_rematch013_inst_rematch013_in_chars,
      rematch013_in_chars_count    => Kernel_rematch013_inst_rematch013_in_chars_count,
      rematch013_in_bus_rreq_valid => Kernel_rematch013_inst_rematch013_in_bus_rreq_valid,
      rematch013_in_bus_rreq_ready => Kernel_rematch013_inst_rematch013_in_bus_rreq_ready,
      rematch013_in_bus_rreq_addr  => Kernel_rematch013_inst_rematch013_in_bus_rreq_addr,
      rematch013_in_bus_rreq_len   => Kernel_rematch013_inst_rematch013_in_bus_rreq_len,
      rematch013_in_bus_rdat_valid => Kernel_rematch013_inst_rematch013_in_bus_rdat_valid,
      rematch013_in_bus_rdat_ready => Kernel_rematch013_inst_rematch013_in_bus_rdat_ready,
      rematch013_in_bus_rdat_data  => Kernel_rematch013_inst_rematch013_in_bus_rdat_data,
      rematch013_in_bus_rdat_last  => Kernel_rematch013_inst_rematch013_in_bus_rdat_last,
      rematch013_in_cmd_valid      => Kernel_rematch013_inst_rematch013_in_cmd_valid,
      rematch013_in_cmd_ready      => Kernel_rematch013_inst_rematch013_in_cmd_ready,
      rematch013_in_cmd_firstIdx   => Kernel_rematch013_inst_rematch013_in_cmd_firstIdx,
      rematch013_in_cmd_lastIdx    => Kernel_rematch013_inst_rematch013_in_cmd_lastIdx,
      rematch013_in_cmd_ctrl       => Kernel_rematch013_inst_rematch013_in_cmd_ctrl,
      rematch013_in_cmd_tag        => Kernel_rematch013_inst_rematch013_in_cmd_tag,
      rematch013_in_unl_valid      => Kernel_rematch013_inst_rematch013_in_unl_valid,
      rematch013_in_unl_ready      => Kernel_rematch013_inst_rematch013_in_unl_ready,
      rematch013_in_unl_tag        => Kernel_rematch013_inst_rematch013_in_unl_tag
    );

  Kernel_rematch014_inst : Kernel_rematch014
    generic map (
      INDEX_WIDTH                      => INDEX_WIDTH,
      TAG_WIDTH                        => TAG_WIDTH,
      REMATCH014_IN_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
      REMATCH014_IN_BUS_DATA_WIDTH     => BUS_DATA_WIDTH,
      REMATCH014_IN_BUS_LEN_WIDTH      => BUS_LEN_WIDTH,
      REMATCH014_IN_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
      REMATCH014_IN_BUS_BURST_MAX_LEN  => BUS_BURST_MAX_LEN
    )
    port map (
      bcd_clk                      => bcd_clk,
      bcd_reset                    => bcd_reset,
      kcd_clk                      => kcd_clk,
      kcd_reset                    => kcd_reset,
      rematch014_in_valid          => Kernel_rematch014_inst_rematch014_in_valid,
      rematch014_in_ready          => Kernel_rematch014_inst_rematch014_in_ready,
      rematch014_in_dvalid         => Kernel_rematch014_inst_rematch014_in_dvalid,
      rematch014_in_last           => Kernel_rematch014_inst_rematch014_in_last,
      rematch014_in_length         => Kernel_rematch014_inst_rematch014_in_length,
      rematch014_in_count          => Kernel_rematch014_inst_rematch014_in_count,
      rematch014_in_chars_valid    => Kernel_rematch014_inst_rematch014_in_chars_valid,
      rematch014_in_chars_ready    => Kernel_rematch014_inst_rematch014_in_chars_ready,
      rematch014_in_chars_dvalid   => Kernel_rematch014_inst_rematch014_in_chars_dvalid,
      rematch014_in_chars_last     => Kernel_rematch014_inst_rematch014_in_chars_last,
      rematch014_in_chars          => Kernel_rematch014_inst_rematch014_in_chars,
      rematch014_in_chars_count    => Kernel_rematch014_inst_rematch014_in_chars_count,
      rematch014_in_bus_rreq_valid => Kernel_rematch014_inst_rematch014_in_bus_rreq_valid,
      rematch014_in_bus_rreq_ready => Kernel_rematch014_inst_rematch014_in_bus_rreq_ready,
      rematch014_in_bus_rreq_addr  => Kernel_rematch014_inst_rematch014_in_bus_rreq_addr,
      rematch014_in_bus_rreq_len   => Kernel_rematch014_inst_rematch014_in_bus_rreq_len,
      rematch014_in_bus_rdat_valid => Kernel_rematch014_inst_rematch014_in_bus_rdat_valid,
      rematch014_in_bus_rdat_ready => Kernel_rematch014_inst_rematch014_in_bus_rdat_ready,
      rematch014_in_bus_rdat_data  => Kernel_rematch014_inst_rematch014_in_bus_rdat_data,
      rematch014_in_bus_rdat_last  => Kernel_rematch014_inst_rematch014_in_bus_rdat_last,
      rematch014_in_cmd_valid      => Kernel_rematch014_inst_rematch014_in_cmd_valid,
      rematch014_in_cmd_ready      => Kernel_rematch014_inst_rematch014_in_cmd_ready,
      rematch014_in_cmd_firstIdx   => Kernel_rematch014_inst_rematch014_in_cmd_firstIdx,
      rematch014_in_cmd_lastIdx    => Kernel_rematch014_inst_rematch014_in_cmd_lastIdx,
      rematch014_in_cmd_ctrl       => Kernel_rematch014_inst_rematch014_in_cmd_ctrl,
      rematch014_in_cmd_tag        => Kernel_rematch014_inst_rematch014_in_cmd_tag,
      rematch014_in_unl_valid      => Kernel_rematch014_inst_rematch014_in_unl_valid,
      rematch014_in_unl_ready      => Kernel_rematch014_inst_rematch014_in_unl_ready,
      rematch014_in_unl_tag        => Kernel_rematch014_inst_rematch014_in_unl_tag
    );

  Kernel_rematch015_inst : Kernel_rematch015
    generic map (
      INDEX_WIDTH                      => INDEX_WIDTH,
      TAG_WIDTH                        => TAG_WIDTH,
      REMATCH015_IN_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
      REMATCH015_IN_BUS_DATA_WIDTH     => BUS_DATA_WIDTH,
      REMATCH015_IN_BUS_LEN_WIDTH      => BUS_LEN_WIDTH,
      REMATCH015_IN_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
      REMATCH015_IN_BUS_BURST_MAX_LEN  => BUS_BURST_MAX_LEN
    )
    port map (
      bcd_clk                      => bcd_clk,
      bcd_reset                    => bcd_reset,
      kcd_clk                      => kcd_clk,
      kcd_reset                    => kcd_reset,
      rematch015_in_valid          => Kernel_rematch015_inst_rematch015_in_valid,
      rematch015_in_ready          => Kernel_rematch015_inst_rematch015_in_ready,
      rematch015_in_dvalid         => Kernel_rematch015_inst_rematch015_in_dvalid,
      rematch015_in_last           => Kernel_rematch015_inst_rematch015_in_last,
      rematch015_in_length         => Kernel_rematch015_inst_rematch015_in_length,
      rematch015_in_count          => Kernel_rematch015_inst_rematch015_in_count,
      rematch015_in_chars_valid    => Kernel_rematch015_inst_rematch015_in_chars_valid,
      rematch015_in_chars_ready    => Kernel_rematch015_inst_rematch015_in_chars_ready,
      rematch015_in_chars_dvalid   => Kernel_rematch015_inst_rematch015_in_chars_dvalid,
      rematch015_in_chars_last     => Kernel_rematch015_inst_rematch015_in_chars_last,
      rematch015_in_chars          => Kernel_rematch015_inst_rematch015_in_chars,
      rematch015_in_chars_count    => Kernel_rematch015_inst_rematch015_in_chars_count,
      rematch015_in_bus_rreq_valid => Kernel_rematch015_inst_rematch015_in_bus_rreq_valid,
      rematch015_in_bus_rreq_ready => Kernel_rematch015_inst_rematch015_in_bus_rreq_ready,
      rematch015_in_bus_rreq_addr  => Kernel_rematch015_inst_rematch015_in_bus_rreq_addr,
      rematch015_in_bus_rreq_len   => Kernel_rematch015_inst_rematch015_in_bus_rreq_len,
      rematch015_in_bus_rdat_valid => Kernel_rematch015_inst_rematch015_in_bus_rdat_valid,
      rematch015_in_bus_rdat_ready => Kernel_rematch015_inst_rematch015_in_bus_rdat_ready,
      rematch015_in_bus_rdat_data  => Kernel_rematch015_inst_rematch015_in_bus_rdat_data,
      rematch015_in_bus_rdat_last  => Kernel_rematch015_inst_rematch015_in_bus_rdat_last,
      rematch015_in_cmd_valid      => Kernel_rematch015_inst_rematch015_in_cmd_valid,
      rematch015_in_cmd_ready      => Kernel_rematch015_inst_rematch015_in_cmd_ready,
      rematch015_in_cmd_firstIdx   => Kernel_rematch015_inst_rematch015_in_cmd_firstIdx,
      rematch015_in_cmd_lastIdx    => Kernel_rematch015_inst_rematch015_in_cmd_lastIdx,
      rematch015_in_cmd_ctrl       => Kernel_rematch015_inst_rematch015_in_cmd_ctrl,
      rematch015_in_cmd_tag        => Kernel_rematch015_inst_rematch015_in_cmd_tag,
      rematch015_in_unl_valid      => Kernel_rematch015_inst_rematch015_in_unl_valid,
      rematch015_in_unl_ready      => Kernel_rematch015_inst_rematch015_in_unl_ready,
      rematch015_in_unl_tag        => Kernel_rematch015_inst_rematch015_in_unl_tag
    );

  RDAW64DW512LW8BS1BM16_inst : BusReadArbiterVec
    generic map (
      BUS_ADDR_WIDTH  => BUS_ADDR_WIDTH,
      BUS_DATA_WIDTH  => BUS_DATA_WIDTH,
      BUS_LEN_WIDTH   => BUS_LEN_WIDTH,
      NUM_SLAVE_PORTS => 16,
      ARB_METHOD      => "RR-STICKY",
      MAX_OUTSTANDING => 4,
      RAM_CONFIG      => "",
      SLV_REQ_SLICES  => true,
      MST_REQ_SLICE   => true,
      MST_DAT_SLICE   => true,
      SLV_DAT_SLICES  => true
    )
    port map (
      bcd_clk        => bcd_clk,
      bcd_reset      => bcd_reset,
      mst_rreq_valid => RDAW64DW512LW8BS1BM16_inst_mst_rreq_valid,
      mst_rreq_ready => RDAW64DW512LW8BS1BM16_inst_mst_rreq_ready,
      mst_rreq_addr  => RDAW64DW512LW8BS1BM16_inst_mst_rreq_addr,
      mst_rreq_len   => RDAW64DW512LW8BS1BM16_inst_mst_rreq_len,
      mst_rdat_valid => RDAW64DW512LW8BS1BM16_inst_mst_rdat_valid,
      mst_rdat_ready => RDAW64DW512LW8BS1BM16_inst_mst_rdat_ready,
      mst_rdat_data  => RDAW64DW512LW8BS1BM16_inst_mst_rdat_data,
      mst_rdat_last  => RDAW64DW512LW8BS1BM16_inst_mst_rdat_last,
      bsv_rreq_valid => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid,
      bsv_rreq_ready => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready,
      bsv_rreq_len   => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len,
      bsv_rreq_addr  => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr,
      bsv_rdat_valid => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid,
      bsv_rdat_ready => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready,
      bsv_rdat_last  => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last,
      bsv_rdat_data  => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data
    );

  rd_mst_rreq_valid                         <= RDAW64DW512LW8BS1BM16_inst_mst_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_mst_rreq_ready <= rd_mst_rreq_ready;
  rd_mst_rreq_addr                          <= RDAW64DW512LW8BS1BM16_inst_mst_rreq_addr;
  rd_mst_rreq_len                           <= RDAW64DW512LW8BS1BM16_inst_mst_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_mst_rdat_valid <= rd_mst_rdat_valid;
  rd_mst_rdat_ready                         <= RDAW64DW512LW8BS1BM16_inst_mst_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_mst_rdat_data  <= rd_mst_rdat_data;
  RDAW64DW512LW8BS1BM16_inst_mst_rdat_last  <= rd_mst_rdat_last;

  Kernel_Nucleus_inst_mmio_awvalid                  <= mmio_awvalid;
  mmio_awready                                      <= Kernel_Nucleus_inst_mmio_awready;
  Kernel_Nucleus_inst_mmio_awaddr                   <= mmio_awaddr;
  Kernel_Nucleus_inst_mmio_wvalid                   <= mmio_wvalid;
  mmio_wready                                       <= Kernel_Nucleus_inst_mmio_wready;
  Kernel_Nucleus_inst_mmio_wdata                    <= mmio_wdata;
  Kernel_Nucleus_inst_mmio_wstrb                    <= mmio_wstrb;
  mmio_bvalid                                       <= Kernel_Nucleus_inst_mmio_bvalid;
  Kernel_Nucleus_inst_mmio_bready                   <= mmio_bready;
  mmio_bresp                                        <= Kernel_Nucleus_inst_mmio_bresp;
  Kernel_Nucleus_inst_mmio_arvalid                  <= mmio_arvalid;
  mmio_arready                                      <= Kernel_Nucleus_inst_mmio_arready;
  Kernel_Nucleus_inst_mmio_araddr                   <= mmio_araddr;
  mmio_rvalid                                       <= Kernel_Nucleus_inst_mmio_rvalid;
  Kernel_Nucleus_inst_mmio_rready                   <= mmio_rready;
  mmio_rdata                                        <= Kernel_Nucleus_inst_mmio_rdata;
  mmio_rresp                                        <= Kernel_Nucleus_inst_mmio_rresp;

  Kernel_Nucleus_inst_rematch000_in_valid           <= Kernel_rematch000_inst_rematch000_in_valid;
  Kernel_rematch000_inst_rematch000_in_ready        <= Kernel_Nucleus_inst_rematch000_in_ready;
  Kernel_Nucleus_inst_rematch000_in_dvalid          <= Kernel_rematch000_inst_rematch000_in_dvalid;
  Kernel_Nucleus_inst_rematch000_in_last            <= Kernel_rematch000_inst_rematch000_in_last;
  Kernel_Nucleus_inst_rematch000_in_length          <= Kernel_rematch000_inst_rematch000_in_length;
  Kernel_Nucleus_inst_rematch000_in_count           <= Kernel_rematch000_inst_rematch000_in_count;
  Kernel_Nucleus_inst_rematch000_in_chars_valid     <= Kernel_rematch000_inst_rematch000_in_chars_valid;
  Kernel_rematch000_inst_rematch000_in_chars_ready  <= Kernel_Nucleus_inst_rematch000_in_chars_ready;
  Kernel_Nucleus_inst_rematch000_in_chars_dvalid    <= Kernel_rematch000_inst_rematch000_in_chars_dvalid;
  Kernel_Nucleus_inst_rematch000_in_chars_last      <= Kernel_rematch000_inst_rematch000_in_chars_last;
  Kernel_Nucleus_inst_rematch000_in_chars           <= Kernel_rematch000_inst_rematch000_in_chars;
  Kernel_Nucleus_inst_rematch000_in_chars_count     <= Kernel_rematch000_inst_rematch000_in_chars_count;

  Kernel_Nucleus_inst_rematch000_in_unl_valid       <= Kernel_rematch000_inst_rematch000_in_unl_valid;
  Kernel_rematch000_inst_rematch000_in_unl_ready    <= Kernel_Nucleus_inst_rematch000_in_unl_ready;
  Kernel_Nucleus_inst_rematch000_in_unl_tag         <= Kernel_rematch000_inst_rematch000_in_unl_tag;

  Kernel_Nucleus_inst_rematch001_in_valid           <= Kernel_rematch001_inst_rematch001_in_valid;
  Kernel_rematch001_inst_rematch001_in_ready        <= Kernel_Nucleus_inst_rematch001_in_ready;
  Kernel_Nucleus_inst_rematch001_in_dvalid          <= Kernel_rematch001_inst_rematch001_in_dvalid;
  Kernel_Nucleus_inst_rematch001_in_last            <= Kernel_rematch001_inst_rematch001_in_last;
  Kernel_Nucleus_inst_rematch001_in_length          <= Kernel_rematch001_inst_rematch001_in_length;
  Kernel_Nucleus_inst_rematch001_in_count           <= Kernel_rematch001_inst_rematch001_in_count;
  Kernel_Nucleus_inst_rematch001_in_chars_valid     <= Kernel_rematch001_inst_rematch001_in_chars_valid;
  Kernel_rematch001_inst_rematch001_in_chars_ready  <= Kernel_Nucleus_inst_rematch001_in_chars_ready;
  Kernel_Nucleus_inst_rematch001_in_chars_dvalid    <= Kernel_rematch001_inst_rematch001_in_chars_dvalid;
  Kernel_Nucleus_inst_rematch001_in_chars_last      <= Kernel_rematch001_inst_rematch001_in_chars_last;
  Kernel_Nucleus_inst_rematch001_in_chars           <= Kernel_rematch001_inst_rematch001_in_chars;
  Kernel_Nucleus_inst_rematch001_in_chars_count     <= Kernel_rematch001_inst_rematch001_in_chars_count;

  Kernel_Nucleus_inst_rematch001_in_unl_valid       <= Kernel_rematch001_inst_rematch001_in_unl_valid;
  Kernel_rematch001_inst_rematch001_in_unl_ready    <= Kernel_Nucleus_inst_rematch001_in_unl_ready;
  Kernel_Nucleus_inst_rematch001_in_unl_tag         <= Kernel_rematch001_inst_rematch001_in_unl_tag;

  Kernel_Nucleus_inst_rematch002_in_valid           <= Kernel_rematch002_inst_rematch002_in_valid;
  Kernel_rematch002_inst_rematch002_in_ready        <= Kernel_Nucleus_inst_rematch002_in_ready;
  Kernel_Nucleus_inst_rematch002_in_dvalid          <= Kernel_rematch002_inst_rematch002_in_dvalid;
  Kernel_Nucleus_inst_rematch002_in_last            <= Kernel_rematch002_inst_rematch002_in_last;
  Kernel_Nucleus_inst_rematch002_in_length          <= Kernel_rematch002_inst_rematch002_in_length;
  Kernel_Nucleus_inst_rematch002_in_count           <= Kernel_rematch002_inst_rematch002_in_count;
  Kernel_Nucleus_inst_rematch002_in_chars_valid     <= Kernel_rematch002_inst_rematch002_in_chars_valid;
  Kernel_rematch002_inst_rematch002_in_chars_ready  <= Kernel_Nucleus_inst_rematch002_in_chars_ready;
  Kernel_Nucleus_inst_rematch002_in_chars_dvalid    <= Kernel_rematch002_inst_rematch002_in_chars_dvalid;
  Kernel_Nucleus_inst_rematch002_in_chars_last      <= Kernel_rematch002_inst_rematch002_in_chars_last;
  Kernel_Nucleus_inst_rematch002_in_chars           <= Kernel_rematch002_inst_rematch002_in_chars;
  Kernel_Nucleus_inst_rematch002_in_chars_count     <= Kernel_rematch002_inst_rematch002_in_chars_count;

  Kernel_Nucleus_inst_rematch002_in_unl_valid       <= Kernel_rematch002_inst_rematch002_in_unl_valid;
  Kernel_rematch002_inst_rematch002_in_unl_ready    <= Kernel_Nucleus_inst_rematch002_in_unl_ready;
  Kernel_Nucleus_inst_rematch002_in_unl_tag         <= Kernel_rematch002_inst_rematch002_in_unl_tag;

  Kernel_Nucleus_inst_rematch003_in_valid           <= Kernel_rematch003_inst_rematch003_in_valid;
  Kernel_rematch003_inst_rematch003_in_ready        <= Kernel_Nucleus_inst_rematch003_in_ready;
  Kernel_Nucleus_inst_rematch003_in_dvalid          <= Kernel_rematch003_inst_rematch003_in_dvalid;
  Kernel_Nucleus_inst_rematch003_in_last            <= Kernel_rematch003_inst_rematch003_in_last;
  Kernel_Nucleus_inst_rematch003_in_length          <= Kernel_rematch003_inst_rematch003_in_length;
  Kernel_Nucleus_inst_rematch003_in_count           <= Kernel_rematch003_inst_rematch003_in_count;
  Kernel_Nucleus_inst_rematch003_in_chars_valid     <= Kernel_rematch003_inst_rematch003_in_chars_valid;
  Kernel_rematch003_inst_rematch003_in_chars_ready  <= Kernel_Nucleus_inst_rematch003_in_chars_ready;
  Kernel_Nucleus_inst_rematch003_in_chars_dvalid    <= Kernel_rematch003_inst_rematch003_in_chars_dvalid;
  Kernel_Nucleus_inst_rematch003_in_chars_last      <= Kernel_rematch003_inst_rematch003_in_chars_last;
  Kernel_Nucleus_inst_rematch003_in_chars           <= Kernel_rematch003_inst_rematch003_in_chars;
  Kernel_Nucleus_inst_rematch003_in_chars_count     <= Kernel_rematch003_inst_rematch003_in_chars_count;

  Kernel_Nucleus_inst_rematch003_in_unl_valid       <= Kernel_rematch003_inst_rematch003_in_unl_valid;
  Kernel_rematch003_inst_rematch003_in_unl_ready    <= Kernel_Nucleus_inst_rematch003_in_unl_ready;
  Kernel_Nucleus_inst_rematch003_in_unl_tag         <= Kernel_rematch003_inst_rematch003_in_unl_tag;

  Kernel_Nucleus_inst_rematch004_in_valid           <= Kernel_rematch004_inst_rematch004_in_valid;
  Kernel_rematch004_inst_rematch004_in_ready        <= Kernel_Nucleus_inst_rematch004_in_ready;
  Kernel_Nucleus_inst_rematch004_in_dvalid          <= Kernel_rematch004_inst_rematch004_in_dvalid;
  Kernel_Nucleus_inst_rematch004_in_last            <= Kernel_rematch004_inst_rematch004_in_last;
  Kernel_Nucleus_inst_rematch004_in_length          <= Kernel_rematch004_inst_rematch004_in_length;
  Kernel_Nucleus_inst_rematch004_in_count           <= Kernel_rematch004_inst_rematch004_in_count;
  Kernel_Nucleus_inst_rematch004_in_chars_valid     <= Kernel_rematch004_inst_rematch004_in_chars_valid;
  Kernel_rematch004_inst_rematch004_in_chars_ready  <= Kernel_Nucleus_inst_rematch004_in_chars_ready;
  Kernel_Nucleus_inst_rematch004_in_chars_dvalid    <= Kernel_rematch004_inst_rematch004_in_chars_dvalid;
  Kernel_Nucleus_inst_rematch004_in_chars_last      <= Kernel_rematch004_inst_rematch004_in_chars_last;
  Kernel_Nucleus_inst_rematch004_in_chars           <= Kernel_rematch004_inst_rematch004_in_chars;
  Kernel_Nucleus_inst_rematch004_in_chars_count     <= Kernel_rematch004_inst_rematch004_in_chars_count;

  Kernel_Nucleus_inst_rematch004_in_unl_valid       <= Kernel_rematch004_inst_rematch004_in_unl_valid;
  Kernel_rematch004_inst_rematch004_in_unl_ready    <= Kernel_Nucleus_inst_rematch004_in_unl_ready;
  Kernel_Nucleus_inst_rematch004_in_unl_tag         <= Kernel_rematch004_inst_rematch004_in_unl_tag;

  Kernel_Nucleus_inst_rematch005_in_valid           <= Kernel_rematch005_inst_rematch005_in_valid;
  Kernel_rematch005_inst_rematch005_in_ready        <= Kernel_Nucleus_inst_rematch005_in_ready;
  Kernel_Nucleus_inst_rematch005_in_dvalid          <= Kernel_rematch005_inst_rematch005_in_dvalid;
  Kernel_Nucleus_inst_rematch005_in_last            <= Kernel_rematch005_inst_rematch005_in_last;
  Kernel_Nucleus_inst_rematch005_in_length          <= Kernel_rematch005_inst_rematch005_in_length;
  Kernel_Nucleus_inst_rematch005_in_count           <= Kernel_rematch005_inst_rematch005_in_count;
  Kernel_Nucleus_inst_rematch005_in_chars_valid     <= Kernel_rematch005_inst_rematch005_in_chars_valid;
  Kernel_rematch005_inst_rematch005_in_chars_ready  <= Kernel_Nucleus_inst_rematch005_in_chars_ready;
  Kernel_Nucleus_inst_rematch005_in_chars_dvalid    <= Kernel_rematch005_inst_rematch005_in_chars_dvalid;
  Kernel_Nucleus_inst_rematch005_in_chars_last      <= Kernel_rematch005_inst_rematch005_in_chars_last;
  Kernel_Nucleus_inst_rematch005_in_chars           <= Kernel_rematch005_inst_rematch005_in_chars;
  Kernel_Nucleus_inst_rematch005_in_chars_count     <= Kernel_rematch005_inst_rematch005_in_chars_count;

  Kernel_Nucleus_inst_rematch005_in_unl_valid       <= Kernel_rematch005_inst_rematch005_in_unl_valid;
  Kernel_rematch005_inst_rematch005_in_unl_ready    <= Kernel_Nucleus_inst_rematch005_in_unl_ready;
  Kernel_Nucleus_inst_rematch005_in_unl_tag         <= Kernel_rematch005_inst_rematch005_in_unl_tag;

  Kernel_Nucleus_inst_rematch006_in_valid           <= Kernel_rematch006_inst_rematch006_in_valid;
  Kernel_rematch006_inst_rematch006_in_ready        <= Kernel_Nucleus_inst_rematch006_in_ready;
  Kernel_Nucleus_inst_rematch006_in_dvalid          <= Kernel_rematch006_inst_rematch006_in_dvalid;
  Kernel_Nucleus_inst_rematch006_in_last            <= Kernel_rematch006_inst_rematch006_in_last;
  Kernel_Nucleus_inst_rematch006_in_length          <= Kernel_rematch006_inst_rematch006_in_length;
  Kernel_Nucleus_inst_rematch006_in_count           <= Kernel_rematch006_inst_rematch006_in_count;
  Kernel_Nucleus_inst_rematch006_in_chars_valid     <= Kernel_rematch006_inst_rematch006_in_chars_valid;
  Kernel_rematch006_inst_rematch006_in_chars_ready  <= Kernel_Nucleus_inst_rematch006_in_chars_ready;
  Kernel_Nucleus_inst_rematch006_in_chars_dvalid    <= Kernel_rematch006_inst_rematch006_in_chars_dvalid;
  Kernel_Nucleus_inst_rematch006_in_chars_last      <= Kernel_rematch006_inst_rematch006_in_chars_last;
  Kernel_Nucleus_inst_rematch006_in_chars           <= Kernel_rematch006_inst_rematch006_in_chars;
  Kernel_Nucleus_inst_rematch006_in_chars_count     <= Kernel_rematch006_inst_rematch006_in_chars_count;

  Kernel_Nucleus_inst_rematch006_in_unl_valid       <= Kernel_rematch006_inst_rematch006_in_unl_valid;
  Kernel_rematch006_inst_rematch006_in_unl_ready    <= Kernel_Nucleus_inst_rematch006_in_unl_ready;
  Kernel_Nucleus_inst_rematch006_in_unl_tag         <= Kernel_rematch006_inst_rematch006_in_unl_tag;

  Kernel_Nucleus_inst_rematch007_in_valid           <= Kernel_rematch007_inst_rematch007_in_valid;
  Kernel_rematch007_inst_rematch007_in_ready        <= Kernel_Nucleus_inst_rematch007_in_ready;
  Kernel_Nucleus_inst_rematch007_in_dvalid          <= Kernel_rematch007_inst_rematch007_in_dvalid;
  Kernel_Nucleus_inst_rematch007_in_last            <= Kernel_rematch007_inst_rematch007_in_last;
  Kernel_Nucleus_inst_rematch007_in_length          <= Kernel_rematch007_inst_rematch007_in_length;
  Kernel_Nucleus_inst_rematch007_in_count           <= Kernel_rematch007_inst_rematch007_in_count;
  Kernel_Nucleus_inst_rematch007_in_chars_valid     <= Kernel_rematch007_inst_rematch007_in_chars_valid;
  Kernel_rematch007_inst_rematch007_in_chars_ready  <= Kernel_Nucleus_inst_rematch007_in_chars_ready;
  Kernel_Nucleus_inst_rematch007_in_chars_dvalid    <= Kernel_rematch007_inst_rematch007_in_chars_dvalid;
  Kernel_Nucleus_inst_rematch007_in_chars_last      <= Kernel_rematch007_inst_rematch007_in_chars_last;
  Kernel_Nucleus_inst_rematch007_in_chars           <= Kernel_rematch007_inst_rematch007_in_chars;
  Kernel_Nucleus_inst_rematch007_in_chars_count     <= Kernel_rematch007_inst_rematch007_in_chars_count;

  Kernel_Nucleus_inst_rematch007_in_unl_valid       <= Kernel_rematch007_inst_rematch007_in_unl_valid;
  Kernel_rematch007_inst_rematch007_in_unl_ready    <= Kernel_Nucleus_inst_rematch007_in_unl_ready;
  Kernel_Nucleus_inst_rematch007_in_unl_tag         <= Kernel_rematch007_inst_rematch007_in_unl_tag;

  Kernel_Nucleus_inst_rematch008_in_valid           <= Kernel_rematch008_inst_rematch008_in_valid;
  Kernel_rematch008_inst_rematch008_in_ready        <= Kernel_Nucleus_inst_rematch008_in_ready;
  Kernel_Nucleus_inst_rematch008_in_dvalid          <= Kernel_rematch008_inst_rematch008_in_dvalid;
  Kernel_Nucleus_inst_rematch008_in_last            <= Kernel_rematch008_inst_rematch008_in_last;
  Kernel_Nucleus_inst_rematch008_in_length          <= Kernel_rematch008_inst_rematch008_in_length;
  Kernel_Nucleus_inst_rematch008_in_count           <= Kernel_rematch008_inst_rematch008_in_count;
  Kernel_Nucleus_inst_rematch008_in_chars_valid     <= Kernel_rematch008_inst_rematch008_in_chars_valid;
  Kernel_rematch008_inst_rematch008_in_chars_ready  <= Kernel_Nucleus_inst_rematch008_in_chars_ready;
  Kernel_Nucleus_inst_rematch008_in_chars_dvalid    <= Kernel_rematch008_inst_rematch008_in_chars_dvalid;
  Kernel_Nucleus_inst_rematch008_in_chars_last      <= Kernel_rematch008_inst_rematch008_in_chars_last;
  Kernel_Nucleus_inst_rematch008_in_chars           <= Kernel_rematch008_inst_rematch008_in_chars;
  Kernel_Nucleus_inst_rematch008_in_chars_count     <= Kernel_rematch008_inst_rematch008_in_chars_count;

  Kernel_Nucleus_inst_rematch008_in_unl_valid       <= Kernel_rematch008_inst_rematch008_in_unl_valid;
  Kernel_rematch008_inst_rematch008_in_unl_ready    <= Kernel_Nucleus_inst_rematch008_in_unl_ready;
  Kernel_Nucleus_inst_rematch008_in_unl_tag         <= Kernel_rematch008_inst_rematch008_in_unl_tag;

  Kernel_Nucleus_inst_rematch009_in_valid           <= Kernel_rematch009_inst_rematch009_in_valid;
  Kernel_rematch009_inst_rematch009_in_ready        <= Kernel_Nucleus_inst_rematch009_in_ready;
  Kernel_Nucleus_inst_rematch009_in_dvalid          <= Kernel_rematch009_inst_rematch009_in_dvalid;
  Kernel_Nucleus_inst_rematch009_in_last            <= Kernel_rematch009_inst_rematch009_in_last;
  Kernel_Nucleus_inst_rematch009_in_length          <= Kernel_rematch009_inst_rematch009_in_length;
  Kernel_Nucleus_inst_rematch009_in_count           <= Kernel_rematch009_inst_rematch009_in_count;
  Kernel_Nucleus_inst_rematch009_in_chars_valid     <= Kernel_rematch009_inst_rematch009_in_chars_valid;
  Kernel_rematch009_inst_rematch009_in_chars_ready  <= Kernel_Nucleus_inst_rematch009_in_chars_ready;
  Kernel_Nucleus_inst_rematch009_in_chars_dvalid    <= Kernel_rematch009_inst_rematch009_in_chars_dvalid;
  Kernel_Nucleus_inst_rematch009_in_chars_last      <= Kernel_rematch009_inst_rematch009_in_chars_last;
  Kernel_Nucleus_inst_rematch009_in_chars           <= Kernel_rematch009_inst_rematch009_in_chars;
  Kernel_Nucleus_inst_rematch009_in_chars_count     <= Kernel_rematch009_inst_rematch009_in_chars_count;

  Kernel_Nucleus_inst_rematch009_in_unl_valid       <= Kernel_rematch009_inst_rematch009_in_unl_valid;
  Kernel_rematch009_inst_rematch009_in_unl_ready    <= Kernel_Nucleus_inst_rematch009_in_unl_ready;
  Kernel_Nucleus_inst_rematch009_in_unl_tag         <= Kernel_rematch009_inst_rematch009_in_unl_tag;

  Kernel_Nucleus_inst_rematch010_in_valid           <= Kernel_rematch010_inst_rematch010_in_valid;
  Kernel_rematch010_inst_rematch010_in_ready        <= Kernel_Nucleus_inst_rematch010_in_ready;
  Kernel_Nucleus_inst_rematch010_in_dvalid          <= Kernel_rematch010_inst_rematch010_in_dvalid;
  Kernel_Nucleus_inst_rematch010_in_last            <= Kernel_rematch010_inst_rematch010_in_last;
  Kernel_Nucleus_inst_rematch010_in_length          <= Kernel_rematch010_inst_rematch010_in_length;
  Kernel_Nucleus_inst_rematch010_in_count           <= Kernel_rematch010_inst_rematch010_in_count;
  Kernel_Nucleus_inst_rematch010_in_chars_valid     <= Kernel_rematch010_inst_rematch010_in_chars_valid;
  Kernel_rematch010_inst_rematch010_in_chars_ready  <= Kernel_Nucleus_inst_rematch010_in_chars_ready;
  Kernel_Nucleus_inst_rematch010_in_chars_dvalid    <= Kernel_rematch010_inst_rematch010_in_chars_dvalid;
  Kernel_Nucleus_inst_rematch010_in_chars_last      <= Kernel_rematch010_inst_rematch010_in_chars_last;
  Kernel_Nucleus_inst_rematch010_in_chars           <= Kernel_rematch010_inst_rematch010_in_chars;
  Kernel_Nucleus_inst_rematch010_in_chars_count     <= Kernel_rematch010_inst_rematch010_in_chars_count;

  Kernel_Nucleus_inst_rematch010_in_unl_valid       <= Kernel_rematch010_inst_rematch010_in_unl_valid;
  Kernel_rematch010_inst_rematch010_in_unl_ready    <= Kernel_Nucleus_inst_rematch010_in_unl_ready;
  Kernel_Nucleus_inst_rematch010_in_unl_tag         <= Kernel_rematch010_inst_rematch010_in_unl_tag;

  Kernel_Nucleus_inst_rematch011_in_valid           <= Kernel_rematch011_inst_rematch011_in_valid;
  Kernel_rematch011_inst_rematch011_in_ready        <= Kernel_Nucleus_inst_rematch011_in_ready;
  Kernel_Nucleus_inst_rematch011_in_dvalid          <= Kernel_rematch011_inst_rematch011_in_dvalid;
  Kernel_Nucleus_inst_rematch011_in_last            <= Kernel_rematch011_inst_rematch011_in_last;
  Kernel_Nucleus_inst_rematch011_in_length          <= Kernel_rematch011_inst_rematch011_in_length;
  Kernel_Nucleus_inst_rematch011_in_count           <= Kernel_rematch011_inst_rematch011_in_count;
  Kernel_Nucleus_inst_rematch011_in_chars_valid     <= Kernel_rematch011_inst_rematch011_in_chars_valid;
  Kernel_rematch011_inst_rematch011_in_chars_ready  <= Kernel_Nucleus_inst_rematch011_in_chars_ready;
  Kernel_Nucleus_inst_rematch011_in_chars_dvalid    <= Kernel_rematch011_inst_rematch011_in_chars_dvalid;
  Kernel_Nucleus_inst_rematch011_in_chars_last      <= Kernel_rematch011_inst_rematch011_in_chars_last;
  Kernel_Nucleus_inst_rematch011_in_chars           <= Kernel_rematch011_inst_rematch011_in_chars;
  Kernel_Nucleus_inst_rematch011_in_chars_count     <= Kernel_rematch011_inst_rematch011_in_chars_count;

  Kernel_Nucleus_inst_rematch011_in_unl_valid       <= Kernel_rematch011_inst_rematch011_in_unl_valid;
  Kernel_rematch011_inst_rematch011_in_unl_ready    <= Kernel_Nucleus_inst_rematch011_in_unl_ready;
  Kernel_Nucleus_inst_rematch011_in_unl_tag         <= Kernel_rematch011_inst_rematch011_in_unl_tag;

  Kernel_Nucleus_inst_rematch012_in_valid           <= Kernel_rematch012_inst_rematch012_in_valid;
  Kernel_rematch012_inst_rematch012_in_ready        <= Kernel_Nucleus_inst_rematch012_in_ready;
  Kernel_Nucleus_inst_rematch012_in_dvalid          <= Kernel_rematch012_inst_rematch012_in_dvalid;
  Kernel_Nucleus_inst_rematch012_in_last            <= Kernel_rematch012_inst_rematch012_in_last;
  Kernel_Nucleus_inst_rematch012_in_length          <= Kernel_rematch012_inst_rematch012_in_length;
  Kernel_Nucleus_inst_rematch012_in_count           <= Kernel_rematch012_inst_rematch012_in_count;
  Kernel_Nucleus_inst_rematch012_in_chars_valid     <= Kernel_rematch012_inst_rematch012_in_chars_valid;
  Kernel_rematch012_inst_rematch012_in_chars_ready  <= Kernel_Nucleus_inst_rematch012_in_chars_ready;
  Kernel_Nucleus_inst_rematch012_in_chars_dvalid    <= Kernel_rematch012_inst_rematch012_in_chars_dvalid;
  Kernel_Nucleus_inst_rematch012_in_chars_last      <= Kernel_rematch012_inst_rematch012_in_chars_last;
  Kernel_Nucleus_inst_rematch012_in_chars           <= Kernel_rematch012_inst_rematch012_in_chars;
  Kernel_Nucleus_inst_rematch012_in_chars_count     <= Kernel_rematch012_inst_rematch012_in_chars_count;

  Kernel_Nucleus_inst_rematch012_in_unl_valid       <= Kernel_rematch012_inst_rematch012_in_unl_valid;
  Kernel_rematch012_inst_rematch012_in_unl_ready    <= Kernel_Nucleus_inst_rematch012_in_unl_ready;
  Kernel_Nucleus_inst_rematch012_in_unl_tag         <= Kernel_rematch012_inst_rematch012_in_unl_tag;

  Kernel_Nucleus_inst_rematch013_in_valid           <= Kernel_rematch013_inst_rematch013_in_valid;
  Kernel_rematch013_inst_rematch013_in_ready        <= Kernel_Nucleus_inst_rematch013_in_ready;
  Kernel_Nucleus_inst_rematch013_in_dvalid          <= Kernel_rematch013_inst_rematch013_in_dvalid;
  Kernel_Nucleus_inst_rematch013_in_last            <= Kernel_rematch013_inst_rematch013_in_last;
  Kernel_Nucleus_inst_rematch013_in_length          <= Kernel_rematch013_inst_rematch013_in_length;
  Kernel_Nucleus_inst_rematch013_in_count           <= Kernel_rematch013_inst_rematch013_in_count;
  Kernel_Nucleus_inst_rematch013_in_chars_valid     <= Kernel_rematch013_inst_rematch013_in_chars_valid;
  Kernel_rematch013_inst_rematch013_in_chars_ready  <= Kernel_Nucleus_inst_rematch013_in_chars_ready;
  Kernel_Nucleus_inst_rematch013_in_chars_dvalid    <= Kernel_rematch013_inst_rematch013_in_chars_dvalid;
  Kernel_Nucleus_inst_rematch013_in_chars_last      <= Kernel_rematch013_inst_rematch013_in_chars_last;
  Kernel_Nucleus_inst_rematch013_in_chars           <= Kernel_rematch013_inst_rematch013_in_chars;
  Kernel_Nucleus_inst_rematch013_in_chars_count     <= Kernel_rematch013_inst_rematch013_in_chars_count;

  Kernel_Nucleus_inst_rematch013_in_unl_valid       <= Kernel_rematch013_inst_rematch013_in_unl_valid;
  Kernel_rematch013_inst_rematch013_in_unl_ready    <= Kernel_Nucleus_inst_rematch013_in_unl_ready;
  Kernel_Nucleus_inst_rematch013_in_unl_tag         <= Kernel_rematch013_inst_rematch013_in_unl_tag;

  Kernel_Nucleus_inst_rematch014_in_valid           <= Kernel_rematch014_inst_rematch014_in_valid;
  Kernel_rematch014_inst_rematch014_in_ready        <= Kernel_Nucleus_inst_rematch014_in_ready;
  Kernel_Nucleus_inst_rematch014_in_dvalid          <= Kernel_rematch014_inst_rematch014_in_dvalid;
  Kernel_Nucleus_inst_rematch014_in_last            <= Kernel_rematch014_inst_rematch014_in_last;
  Kernel_Nucleus_inst_rematch014_in_length          <= Kernel_rematch014_inst_rematch014_in_length;
  Kernel_Nucleus_inst_rematch014_in_count           <= Kernel_rematch014_inst_rematch014_in_count;
  Kernel_Nucleus_inst_rematch014_in_chars_valid     <= Kernel_rematch014_inst_rematch014_in_chars_valid;
  Kernel_rematch014_inst_rematch014_in_chars_ready  <= Kernel_Nucleus_inst_rematch014_in_chars_ready;
  Kernel_Nucleus_inst_rematch014_in_chars_dvalid    <= Kernel_rematch014_inst_rematch014_in_chars_dvalid;
  Kernel_Nucleus_inst_rematch014_in_chars_last      <= Kernel_rematch014_inst_rematch014_in_chars_last;
  Kernel_Nucleus_inst_rematch014_in_chars           <= Kernel_rematch014_inst_rematch014_in_chars;
  Kernel_Nucleus_inst_rematch014_in_chars_count     <= Kernel_rematch014_inst_rematch014_in_chars_count;

  Kernel_Nucleus_inst_rematch014_in_unl_valid       <= Kernel_rematch014_inst_rematch014_in_unl_valid;
  Kernel_rematch014_inst_rematch014_in_unl_ready    <= Kernel_Nucleus_inst_rematch014_in_unl_ready;
  Kernel_Nucleus_inst_rematch014_in_unl_tag         <= Kernel_rematch014_inst_rematch014_in_unl_tag;

  Kernel_Nucleus_inst_rematch015_in_valid           <= Kernel_rematch015_inst_rematch015_in_valid;
  Kernel_rematch015_inst_rematch015_in_ready        <= Kernel_Nucleus_inst_rematch015_in_ready;
  Kernel_Nucleus_inst_rematch015_in_dvalid          <= Kernel_rematch015_inst_rematch015_in_dvalid;
  Kernel_Nucleus_inst_rematch015_in_last            <= Kernel_rematch015_inst_rematch015_in_last;
  Kernel_Nucleus_inst_rematch015_in_length          <= Kernel_rematch015_inst_rematch015_in_length;
  Kernel_Nucleus_inst_rematch015_in_count           <= Kernel_rematch015_inst_rematch015_in_count;
  Kernel_Nucleus_inst_rematch015_in_chars_valid     <= Kernel_rematch015_inst_rematch015_in_chars_valid;
  Kernel_rematch015_inst_rematch015_in_chars_ready  <= Kernel_Nucleus_inst_rematch015_in_chars_ready;
  Kernel_Nucleus_inst_rematch015_in_chars_dvalid    <= Kernel_rematch015_inst_rematch015_in_chars_dvalid;
  Kernel_Nucleus_inst_rematch015_in_chars_last      <= Kernel_rematch015_inst_rematch015_in_chars_last;
  Kernel_Nucleus_inst_rematch015_in_chars           <= Kernel_rematch015_inst_rematch015_in_chars;
  Kernel_Nucleus_inst_rematch015_in_chars_count     <= Kernel_rematch015_inst_rematch015_in_chars_count;

  Kernel_Nucleus_inst_rematch015_in_unl_valid       <= Kernel_rematch015_inst_rematch015_in_unl_valid;
  Kernel_rematch015_inst_rematch015_in_unl_ready    <= Kernel_Nucleus_inst_rematch015_in_unl_ready;
  Kernel_Nucleus_inst_rematch015_in_unl_tag         <= Kernel_rematch015_inst_rematch015_in_unl_tag;

  Kernel_rematch000_inst_rematch000_in_cmd_valid    <= Kernel_Nucleus_inst_rematch000_in_cmd_valid;
  Kernel_Nucleus_inst_rematch000_in_cmd_ready       <= Kernel_rematch000_inst_rematch000_in_cmd_ready;
  Kernel_rematch000_inst_rematch000_in_cmd_firstIdx <= Kernel_Nucleus_inst_rematch000_in_cmd_firstIdx;
  Kernel_rematch000_inst_rematch000_in_cmd_lastIdx  <= Kernel_Nucleus_inst_rematch000_in_cmd_lastIdx;
  Kernel_rematch000_inst_rematch000_in_cmd_ctrl     <= Kernel_Nucleus_inst_rematch000_in_cmd_ctrl;
  Kernel_rematch000_inst_rematch000_in_cmd_tag      <= Kernel_Nucleus_inst_rematch000_in_cmd_tag;

  Kernel_rematch001_inst_rematch001_in_cmd_valid    <= Kernel_Nucleus_inst_rematch001_in_cmd_valid;
  Kernel_Nucleus_inst_rematch001_in_cmd_ready       <= Kernel_rematch001_inst_rematch001_in_cmd_ready;
  Kernel_rematch001_inst_rematch001_in_cmd_firstIdx <= Kernel_Nucleus_inst_rematch001_in_cmd_firstIdx;
  Kernel_rematch001_inst_rematch001_in_cmd_lastIdx  <= Kernel_Nucleus_inst_rematch001_in_cmd_lastIdx;
  Kernel_rematch001_inst_rematch001_in_cmd_ctrl     <= Kernel_Nucleus_inst_rematch001_in_cmd_ctrl;
  Kernel_rematch001_inst_rematch001_in_cmd_tag      <= Kernel_Nucleus_inst_rematch001_in_cmd_tag;

  Kernel_rematch002_inst_rematch002_in_cmd_valid    <= Kernel_Nucleus_inst_rematch002_in_cmd_valid;
  Kernel_Nucleus_inst_rematch002_in_cmd_ready       <= Kernel_rematch002_inst_rematch002_in_cmd_ready;
  Kernel_rematch002_inst_rematch002_in_cmd_firstIdx <= Kernel_Nucleus_inst_rematch002_in_cmd_firstIdx;
  Kernel_rematch002_inst_rematch002_in_cmd_lastIdx  <= Kernel_Nucleus_inst_rematch002_in_cmd_lastIdx;
  Kernel_rematch002_inst_rematch002_in_cmd_ctrl     <= Kernel_Nucleus_inst_rematch002_in_cmd_ctrl;
  Kernel_rematch002_inst_rematch002_in_cmd_tag      <= Kernel_Nucleus_inst_rematch002_in_cmd_tag;

  Kernel_rematch003_inst_rematch003_in_cmd_valid    <= Kernel_Nucleus_inst_rematch003_in_cmd_valid;
  Kernel_Nucleus_inst_rematch003_in_cmd_ready       <= Kernel_rematch003_inst_rematch003_in_cmd_ready;
  Kernel_rematch003_inst_rematch003_in_cmd_firstIdx <= Kernel_Nucleus_inst_rematch003_in_cmd_firstIdx;
  Kernel_rematch003_inst_rematch003_in_cmd_lastIdx  <= Kernel_Nucleus_inst_rematch003_in_cmd_lastIdx;
  Kernel_rematch003_inst_rematch003_in_cmd_ctrl     <= Kernel_Nucleus_inst_rematch003_in_cmd_ctrl;
  Kernel_rematch003_inst_rematch003_in_cmd_tag      <= Kernel_Nucleus_inst_rematch003_in_cmd_tag;

  Kernel_rematch004_inst_rematch004_in_cmd_valid    <= Kernel_Nucleus_inst_rematch004_in_cmd_valid;
  Kernel_Nucleus_inst_rematch004_in_cmd_ready       <= Kernel_rematch004_inst_rematch004_in_cmd_ready;
  Kernel_rematch004_inst_rematch004_in_cmd_firstIdx <= Kernel_Nucleus_inst_rematch004_in_cmd_firstIdx;
  Kernel_rematch004_inst_rematch004_in_cmd_lastIdx  <= Kernel_Nucleus_inst_rematch004_in_cmd_lastIdx;
  Kernel_rematch004_inst_rematch004_in_cmd_ctrl     <= Kernel_Nucleus_inst_rematch004_in_cmd_ctrl;
  Kernel_rematch004_inst_rematch004_in_cmd_tag      <= Kernel_Nucleus_inst_rematch004_in_cmd_tag;

  Kernel_rematch005_inst_rematch005_in_cmd_valid    <= Kernel_Nucleus_inst_rematch005_in_cmd_valid;
  Kernel_Nucleus_inst_rematch005_in_cmd_ready       <= Kernel_rematch005_inst_rematch005_in_cmd_ready;
  Kernel_rematch005_inst_rematch005_in_cmd_firstIdx <= Kernel_Nucleus_inst_rematch005_in_cmd_firstIdx;
  Kernel_rematch005_inst_rematch005_in_cmd_lastIdx  <= Kernel_Nucleus_inst_rematch005_in_cmd_lastIdx;
  Kernel_rematch005_inst_rematch005_in_cmd_ctrl     <= Kernel_Nucleus_inst_rematch005_in_cmd_ctrl;
  Kernel_rematch005_inst_rematch005_in_cmd_tag      <= Kernel_Nucleus_inst_rematch005_in_cmd_tag;

  Kernel_rematch006_inst_rematch006_in_cmd_valid    <= Kernel_Nucleus_inst_rematch006_in_cmd_valid;
  Kernel_Nucleus_inst_rematch006_in_cmd_ready       <= Kernel_rematch006_inst_rematch006_in_cmd_ready;
  Kernel_rematch006_inst_rematch006_in_cmd_firstIdx <= Kernel_Nucleus_inst_rematch006_in_cmd_firstIdx;
  Kernel_rematch006_inst_rematch006_in_cmd_lastIdx  <= Kernel_Nucleus_inst_rematch006_in_cmd_lastIdx;
  Kernel_rematch006_inst_rematch006_in_cmd_ctrl     <= Kernel_Nucleus_inst_rematch006_in_cmd_ctrl;
  Kernel_rematch006_inst_rematch006_in_cmd_tag      <= Kernel_Nucleus_inst_rematch006_in_cmd_tag;

  Kernel_rematch007_inst_rematch007_in_cmd_valid    <= Kernel_Nucleus_inst_rematch007_in_cmd_valid;
  Kernel_Nucleus_inst_rematch007_in_cmd_ready       <= Kernel_rematch007_inst_rematch007_in_cmd_ready;
  Kernel_rematch007_inst_rematch007_in_cmd_firstIdx <= Kernel_Nucleus_inst_rematch007_in_cmd_firstIdx;
  Kernel_rematch007_inst_rematch007_in_cmd_lastIdx  <= Kernel_Nucleus_inst_rematch007_in_cmd_lastIdx;
  Kernel_rematch007_inst_rematch007_in_cmd_ctrl     <= Kernel_Nucleus_inst_rematch007_in_cmd_ctrl;
  Kernel_rematch007_inst_rematch007_in_cmd_tag      <= Kernel_Nucleus_inst_rematch007_in_cmd_tag;

  Kernel_rematch008_inst_rematch008_in_cmd_valid    <= Kernel_Nucleus_inst_rematch008_in_cmd_valid;
  Kernel_Nucleus_inst_rematch008_in_cmd_ready       <= Kernel_rematch008_inst_rematch008_in_cmd_ready;
  Kernel_rematch008_inst_rematch008_in_cmd_firstIdx <= Kernel_Nucleus_inst_rematch008_in_cmd_firstIdx;
  Kernel_rematch008_inst_rematch008_in_cmd_lastIdx  <= Kernel_Nucleus_inst_rematch008_in_cmd_lastIdx;
  Kernel_rematch008_inst_rematch008_in_cmd_ctrl     <= Kernel_Nucleus_inst_rematch008_in_cmd_ctrl;
  Kernel_rematch008_inst_rematch008_in_cmd_tag      <= Kernel_Nucleus_inst_rematch008_in_cmd_tag;

  Kernel_rematch009_inst_rematch009_in_cmd_valid    <= Kernel_Nucleus_inst_rematch009_in_cmd_valid;
  Kernel_Nucleus_inst_rematch009_in_cmd_ready       <= Kernel_rematch009_inst_rematch009_in_cmd_ready;
  Kernel_rematch009_inst_rematch009_in_cmd_firstIdx <= Kernel_Nucleus_inst_rematch009_in_cmd_firstIdx;
  Kernel_rematch009_inst_rematch009_in_cmd_lastIdx  <= Kernel_Nucleus_inst_rematch009_in_cmd_lastIdx;
  Kernel_rematch009_inst_rematch009_in_cmd_ctrl     <= Kernel_Nucleus_inst_rematch009_in_cmd_ctrl;
  Kernel_rematch009_inst_rematch009_in_cmd_tag      <= Kernel_Nucleus_inst_rematch009_in_cmd_tag;

  Kernel_rematch010_inst_rematch010_in_cmd_valid    <= Kernel_Nucleus_inst_rematch010_in_cmd_valid;
  Kernel_Nucleus_inst_rematch010_in_cmd_ready       <= Kernel_rematch010_inst_rematch010_in_cmd_ready;
  Kernel_rematch010_inst_rematch010_in_cmd_firstIdx <= Kernel_Nucleus_inst_rematch010_in_cmd_firstIdx;
  Kernel_rematch010_inst_rematch010_in_cmd_lastIdx  <= Kernel_Nucleus_inst_rematch010_in_cmd_lastIdx;
  Kernel_rematch010_inst_rematch010_in_cmd_ctrl     <= Kernel_Nucleus_inst_rematch010_in_cmd_ctrl;
  Kernel_rematch010_inst_rematch010_in_cmd_tag      <= Kernel_Nucleus_inst_rematch010_in_cmd_tag;

  Kernel_rematch011_inst_rematch011_in_cmd_valid    <= Kernel_Nucleus_inst_rematch011_in_cmd_valid;
  Kernel_Nucleus_inst_rematch011_in_cmd_ready       <= Kernel_rematch011_inst_rematch011_in_cmd_ready;
  Kernel_rematch011_inst_rematch011_in_cmd_firstIdx <= Kernel_Nucleus_inst_rematch011_in_cmd_firstIdx;
  Kernel_rematch011_inst_rematch011_in_cmd_lastIdx  <= Kernel_Nucleus_inst_rematch011_in_cmd_lastIdx;
  Kernel_rematch011_inst_rematch011_in_cmd_ctrl     <= Kernel_Nucleus_inst_rematch011_in_cmd_ctrl;
  Kernel_rematch011_inst_rematch011_in_cmd_tag      <= Kernel_Nucleus_inst_rematch011_in_cmd_tag;

  Kernel_rematch012_inst_rematch012_in_cmd_valid    <= Kernel_Nucleus_inst_rematch012_in_cmd_valid;
  Kernel_Nucleus_inst_rematch012_in_cmd_ready       <= Kernel_rematch012_inst_rematch012_in_cmd_ready;
  Kernel_rematch012_inst_rematch012_in_cmd_firstIdx <= Kernel_Nucleus_inst_rematch012_in_cmd_firstIdx;
  Kernel_rematch012_inst_rematch012_in_cmd_lastIdx  <= Kernel_Nucleus_inst_rematch012_in_cmd_lastIdx;
  Kernel_rematch012_inst_rematch012_in_cmd_ctrl     <= Kernel_Nucleus_inst_rematch012_in_cmd_ctrl;
  Kernel_rematch012_inst_rematch012_in_cmd_tag      <= Kernel_Nucleus_inst_rematch012_in_cmd_tag;

  Kernel_rematch013_inst_rematch013_in_cmd_valid    <= Kernel_Nucleus_inst_rematch013_in_cmd_valid;
  Kernel_Nucleus_inst_rematch013_in_cmd_ready       <= Kernel_rematch013_inst_rematch013_in_cmd_ready;
  Kernel_rematch013_inst_rematch013_in_cmd_firstIdx <= Kernel_Nucleus_inst_rematch013_in_cmd_firstIdx;
  Kernel_rematch013_inst_rematch013_in_cmd_lastIdx  <= Kernel_Nucleus_inst_rematch013_in_cmd_lastIdx;
  Kernel_rematch013_inst_rematch013_in_cmd_ctrl     <= Kernel_Nucleus_inst_rematch013_in_cmd_ctrl;
  Kernel_rematch013_inst_rematch013_in_cmd_tag      <= Kernel_Nucleus_inst_rematch013_in_cmd_tag;

  Kernel_rematch014_inst_rematch014_in_cmd_valid    <= Kernel_Nucleus_inst_rematch014_in_cmd_valid;
  Kernel_Nucleus_inst_rematch014_in_cmd_ready       <= Kernel_rematch014_inst_rematch014_in_cmd_ready;
  Kernel_rematch014_inst_rematch014_in_cmd_firstIdx <= Kernel_Nucleus_inst_rematch014_in_cmd_firstIdx;
  Kernel_rematch014_inst_rematch014_in_cmd_lastIdx  <= Kernel_Nucleus_inst_rematch014_in_cmd_lastIdx;
  Kernel_rematch014_inst_rematch014_in_cmd_ctrl     <= Kernel_Nucleus_inst_rematch014_in_cmd_ctrl;
  Kernel_rematch014_inst_rematch014_in_cmd_tag      <= Kernel_Nucleus_inst_rematch014_in_cmd_tag;

  Kernel_rematch015_inst_rematch015_in_cmd_valid    <= Kernel_Nucleus_inst_rematch015_in_cmd_valid;
  Kernel_Nucleus_inst_rematch015_in_cmd_ready       <= Kernel_rematch015_inst_rematch015_in_cmd_ready;
  Kernel_rematch015_inst_rematch015_in_cmd_firstIdx <= Kernel_Nucleus_inst_rematch015_in_cmd_firstIdx;
  Kernel_rematch015_inst_rematch015_in_cmd_lastIdx  <= Kernel_Nucleus_inst_rematch015_in_cmd_lastIdx;
  Kernel_rematch015_inst_rematch015_in_cmd_ctrl     <= Kernel_Nucleus_inst_rematch015_in_cmd_ctrl;
  Kernel_rematch015_inst_rematch015_in_cmd_tag      <= Kernel_Nucleus_inst_rematch015_in_cmd_tag;

  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(0)                                                          <= Kernel_rematch000_inst_rematch000_in_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(1)                                                          <= Kernel_rematch001_inst_rematch001_in_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(2)                                                          <= Kernel_rematch002_inst_rematch002_in_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(3)                                                          <= Kernel_rematch003_inst_rematch003_in_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(4)                                                          <= Kernel_rematch004_inst_rematch004_in_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(5)                                                          <= Kernel_rematch005_inst_rematch005_in_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(6)                                                          <= Kernel_rematch006_inst_rematch006_in_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(7)                                                          <= Kernel_rematch007_inst_rematch007_in_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(8)                                                          <= Kernel_rematch008_inst_rematch008_in_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(9)                                                          <= Kernel_rematch009_inst_rematch009_in_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(10)                                                         <= Kernel_rematch010_inst_rematch010_in_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(11)                                                         <= Kernel_rematch011_inst_rematch011_in_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(12)                                                         <= Kernel_rematch012_inst_rematch012_in_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(13)                                                         <= Kernel_rematch013_inst_rematch013_in_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(14)                                                         <= Kernel_rematch014_inst_rematch014_in_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(15)                                                         <= Kernel_rematch015_inst_rematch015_in_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH-1 downto 0)                                     <= Kernel_rematch000_inst_rematch000_in_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH)           <= Kernel_rematch001_inst_rematch001_in_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH*2+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*2)       <= Kernel_rematch002_inst_rematch002_in_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH*3+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*3)       <= Kernel_rematch003_inst_rematch003_in_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH*4+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*4)       <= Kernel_rematch004_inst_rematch004_in_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH*5+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*5)       <= Kernel_rematch005_inst_rematch005_in_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH*6+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*6)       <= Kernel_rematch006_inst_rematch006_in_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH*7+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*7)       <= Kernel_rematch007_inst_rematch007_in_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH*8+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*8)       <= Kernel_rematch008_inst_rematch008_in_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH*9+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*9)       <= Kernel_rematch009_inst_rematch009_in_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH*10+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*10)     <= Kernel_rematch010_inst_rematch010_in_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH*11+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*11)     <= Kernel_rematch011_inst_rematch011_in_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH*12+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*12)     <= Kernel_rematch012_inst_rematch012_in_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH*13+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*13)     <= Kernel_rematch013_inst_rematch013_in_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH*14+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*14)     <= Kernel_rematch014_inst_rematch014_in_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH*15+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*15)     <= Kernel_rematch015_inst_rematch015_in_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH-1 downto 0)                                   <= Kernel_rematch000_inst_rematch000_in_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH)       <= Kernel_rematch001_inst_rematch001_in_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH*2+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*2)   <= Kernel_rematch002_inst_rematch002_in_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH*3+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*3)   <= Kernel_rematch003_inst_rematch003_in_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH*4+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*4)   <= Kernel_rematch004_inst_rematch004_in_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH*5+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*5)   <= Kernel_rematch005_inst_rematch005_in_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH*6+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*6)   <= Kernel_rematch006_inst_rematch006_in_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH*7+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*7)   <= Kernel_rematch007_inst_rematch007_in_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH*8+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*8)   <= Kernel_rematch008_inst_rematch008_in_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH*9+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*9)   <= Kernel_rematch009_inst_rematch009_in_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH*10+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*10) <= Kernel_rematch010_inst_rematch010_in_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH*11+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*11) <= Kernel_rematch011_inst_rematch011_in_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH*12+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*12) <= Kernel_rematch012_inst_rematch012_in_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH*13+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*13) <= Kernel_rematch013_inst_rematch013_in_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH*14+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*14) <= Kernel_rematch014_inst_rematch014_in_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH*15+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*15) <= Kernel_rematch015_inst_rematch015_in_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(0)                                                          <= Kernel_rematch000_inst_rematch000_in_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(1)                                                          <= Kernel_rematch001_inst_rematch001_in_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(2)                                                          <= Kernel_rematch002_inst_rematch002_in_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(3)                                                          <= Kernel_rematch003_inst_rematch003_in_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(4)                                                          <= Kernel_rematch004_inst_rematch004_in_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(5)                                                          <= Kernel_rematch005_inst_rematch005_in_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(6)                                                          <= Kernel_rematch006_inst_rematch006_in_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(7)                                                          <= Kernel_rematch007_inst_rematch007_in_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(8)                                                          <= Kernel_rematch008_inst_rematch008_in_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(9)                                                          <= Kernel_rematch009_inst_rematch009_in_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(10)                                                         <= Kernel_rematch010_inst_rematch010_in_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(11)                                                         <= Kernel_rematch011_inst_rematch011_in_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(12)                                                         <= Kernel_rematch012_inst_rematch012_in_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(13)                                                         <= Kernel_rematch013_inst_rematch013_in_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(14)                                                         <= Kernel_rematch014_inst_rematch014_in_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(15)                                                         <= Kernel_rematch015_inst_rematch015_in_bus_rdat_ready;
  Kernel_rematch015_inst_rematch015_in_bus_rreq_ready                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(15);
  Kernel_rematch015_inst_rematch015_in_bus_rdat_valid                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(15);
  Kernel_rematch015_inst_rematch015_in_bus_rdat_last                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(15);
  Kernel_rematch015_inst_rematch015_in_bus_rdat_data                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH*15+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*15);
  Kernel_rematch014_inst_rematch014_in_bus_rreq_ready                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(14);
  Kernel_rematch014_inst_rematch014_in_bus_rdat_valid                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(14);
  Kernel_rematch014_inst_rematch014_in_bus_rdat_last                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(14);
  Kernel_rematch014_inst_rematch014_in_bus_rdat_data                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH*14+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*14);
  Kernel_rematch013_inst_rematch013_in_bus_rreq_ready                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(13);
  Kernel_rematch013_inst_rematch013_in_bus_rdat_valid                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(13);
  Kernel_rematch013_inst_rematch013_in_bus_rdat_last                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(13);
  Kernel_rematch013_inst_rematch013_in_bus_rdat_data                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH*13+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*13);
  Kernel_rematch012_inst_rematch012_in_bus_rreq_ready                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(12);
  Kernel_rematch012_inst_rematch012_in_bus_rdat_valid                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(12);
  Kernel_rematch012_inst_rematch012_in_bus_rdat_last                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(12);
  Kernel_rematch012_inst_rematch012_in_bus_rdat_data                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH*12+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*12);
  Kernel_rematch011_inst_rematch011_in_bus_rreq_ready                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(11);
  Kernel_rematch011_inst_rematch011_in_bus_rdat_valid                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(11);
  Kernel_rematch011_inst_rematch011_in_bus_rdat_last                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(11);
  Kernel_rematch011_inst_rematch011_in_bus_rdat_data                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH*11+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*11);
  Kernel_rematch010_inst_rematch010_in_bus_rreq_ready                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(10);
  Kernel_rematch010_inst_rematch010_in_bus_rdat_valid                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(10);
  Kernel_rematch010_inst_rematch010_in_bus_rdat_last                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(10);
  Kernel_rematch010_inst_rematch010_in_bus_rdat_data                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH*10+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*10);
  Kernel_rematch009_inst_rematch009_in_bus_rreq_ready                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(9);
  Kernel_rematch009_inst_rematch009_in_bus_rdat_valid                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(9);
  Kernel_rematch009_inst_rematch009_in_bus_rdat_last                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(9);
  Kernel_rematch009_inst_rematch009_in_bus_rdat_data                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH*9+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*9);
  Kernel_rematch008_inst_rematch008_in_bus_rreq_ready                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(8);
  Kernel_rematch008_inst_rematch008_in_bus_rdat_valid                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(8);
  Kernel_rematch008_inst_rematch008_in_bus_rdat_last                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(8);
  Kernel_rematch008_inst_rematch008_in_bus_rdat_data                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH*8+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*8);
  Kernel_rematch007_inst_rematch007_in_bus_rreq_ready                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(7);
  Kernel_rematch007_inst_rematch007_in_bus_rdat_valid                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(7);
  Kernel_rematch007_inst_rematch007_in_bus_rdat_last                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(7);
  Kernel_rematch007_inst_rematch007_in_bus_rdat_data                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH*7+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*7);
  Kernel_rematch006_inst_rematch006_in_bus_rreq_ready                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(6);
  Kernel_rematch006_inst_rematch006_in_bus_rdat_valid                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(6);
  Kernel_rematch006_inst_rematch006_in_bus_rdat_last                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(6);
  Kernel_rematch006_inst_rematch006_in_bus_rdat_data                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH*6+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*6);
  Kernel_rematch005_inst_rematch005_in_bus_rreq_ready                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(5);
  Kernel_rematch005_inst_rematch005_in_bus_rdat_valid                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(5);
  Kernel_rematch005_inst_rematch005_in_bus_rdat_last                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(5);
  Kernel_rematch005_inst_rematch005_in_bus_rdat_data                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH*5+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*5);
  Kernel_rematch004_inst_rematch004_in_bus_rreq_ready                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(4);
  Kernel_rematch004_inst_rematch004_in_bus_rdat_valid                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(4);
  Kernel_rematch004_inst_rematch004_in_bus_rdat_last                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(4);
  Kernel_rematch004_inst_rematch004_in_bus_rdat_data                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH*4+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*4);
  Kernel_rematch003_inst_rematch003_in_bus_rreq_ready                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(3);
  Kernel_rematch003_inst_rematch003_in_bus_rdat_valid                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(3);
  Kernel_rematch003_inst_rematch003_in_bus_rdat_last                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(3);
  Kernel_rematch003_inst_rematch003_in_bus_rdat_data                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH*3+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*3);
  Kernel_rematch002_inst_rematch002_in_bus_rreq_ready                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(2);
  Kernel_rematch002_inst_rematch002_in_bus_rdat_valid                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(2);
  Kernel_rematch002_inst_rematch002_in_bus_rdat_last                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(2);
  Kernel_rematch002_inst_rematch002_in_bus_rdat_data                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH*2+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*2);
  Kernel_rematch001_inst_rematch001_in_bus_rreq_ready                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(1);
  Kernel_rematch001_inst_rematch001_in_bus_rdat_valid                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(1);
  Kernel_rematch001_inst_rematch001_in_bus_rdat_last                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(1);
  Kernel_rematch001_inst_rematch001_in_bus_rdat_data                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH);
  Kernel_rematch000_inst_rematch000_in_bus_rreq_ready                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(0);
  Kernel_rematch000_inst_rematch000_in_bus_rdat_valid                                                   <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(0);
  Kernel_rematch000_inst_rematch000_in_bus_rdat_last                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(0);
  Kernel_rematch000_inst_rematch000_in_bus_rdat_data                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH-1 downto 0);

end architecture;
